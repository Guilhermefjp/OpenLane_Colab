magic
tech sky130A
magscale 1 2
timestamp 1571791925
<< checkpaint >>
rect -3932 -3924 23239 25140
<< metal1 >>
rect 1104 18992 18124 19088
rect 2148 18680 2176 18748
rect 4356 18680 4384 18748
rect 4540 18720 4844 18748
rect 7484 18720 10456 18748
rect 2148 18652 3832 18680
rect 4356 18652 4752 18680
rect 4172 18584 4660 18612
rect 10428 18584 10548 18612
rect 1104 18448 18124 18544
rect 5460 18380 5948 18408
rect 6012 18340 6040 18408
rect 2516 18312 3648 18340
rect 4554 18312 5120 18340
rect 5552 18312 6040 18340
rect 1964 18244 2084 18272
rect 2516 18244 2544 18312
rect 5184 18204 5212 18272
rect 5736 18244 5856 18272
rect 6564 18244 7512 18272
rect 6564 18204 6592 18244
rect 2884 18176 3004 18204
rect 3068 18176 3188 18204
rect 5184 18176 6592 18204
rect 9048 18176 9444 18204
rect 3160 18040 3188 18176
rect 7300 18040 7788 18068
rect 1104 17904 18124 18000
rect 1504 17836 2820 17864
rect 3160 17836 3280 17864
rect 3252 17796 3280 17836
rect 3252 17768 5120 17796
rect 8772 17768 8984 17796
rect 10336 17768 12204 17796
rect 3252 17728 3280 17768
rect 5092 17728 5120 17768
rect 1780 17700 3280 17728
rect 3620 17700 3832 17728
rect 5092 17700 6684 17728
rect 8418 17632 8524 17660
rect 10336 17592 10364 17768
rect 10428 17700 12020 17728
rect 1596 17564 1794 17592
rect 5368 17564 5672 17592
rect 8772 17564 9168 17592
rect 9876 17524 9904 17592
rect 10336 17564 10732 17592
rect 10888 17524 10916 17660
rect 11256 17632 11376 17660
rect 12176 17632 12204 17768
rect 6104 17496 6868 17524
rect 9876 17496 10916 17524
rect 11808 17496 11928 17524
rect 11992 17496 12388 17524
rect 1104 17360 18124 17456
rect 2240 17292 3740 17320
rect 3344 17224 3464 17252
rect 3804 17184 3832 17320
rect 3988 17224 4660 17252
rect 5368 17224 5672 17252
rect 2976 17156 3832 17184
rect 8496 17184 8524 17320
rect 9048 17292 9536 17320
rect 9692 17224 10364 17252
rect 8496 17156 8892 17184
rect 9324 17156 9444 17184
rect 9416 17116 9444 17156
rect 10704 17116 10732 17320
rect 10888 17292 12020 17320
rect 10888 17224 10916 17292
rect 10796 17156 11008 17184
rect 11164 17116 11192 17184
rect 6656 17088 6776 17116
rect 7668 17088 8708 17116
rect 9232 17088 11192 17116
rect 11348 17088 11560 17116
rect 9232 16980 9260 17088
rect 7116 16952 9260 16980
rect 11164 16980 11192 17088
rect 11164 16952 11836 16980
rect 13096 16952 13308 16980
rect 1104 16816 18124 16912
rect 10704 16748 10916 16776
rect 12544 16748 12664 16776
rect 3804 16680 7144 16708
rect 1412 16612 1808 16640
rect 2884 16612 4384 16640
rect 4356 16574 4384 16612
rect 3804 16436 3832 16572
rect 4356 16546 4421 16574
rect 4356 16544 4384 16546
rect 4540 16544 4568 16680
rect 4632 16612 5488 16640
rect 5368 16572 5396 16612
rect 5331 16544 5396 16572
rect 5552 16544 5580 16680
rect 5644 16612 6040 16640
rect 6932 16612 7052 16640
rect 7116 16572 7144 16680
rect 10428 16680 11376 16708
rect 10428 16640 10456 16680
rect 9140 16612 10456 16640
rect 12544 16612 14320 16640
rect 12544 16572 12572 16612
rect 5736 16544 6132 16572
rect 7116 16544 7420 16572
rect 7576 16544 7696 16572
rect 10796 16544 12572 16572
rect 4632 16476 4752 16504
rect 3160 16408 3832 16436
rect 1104 16272 18124 16368
rect 2884 16204 3004 16232
rect 3068 16204 4200 16232
rect 6012 16204 6132 16232
rect 6196 16204 6500 16232
rect 9416 16204 9628 16232
rect 10152 16204 10272 16232
rect 1688 16136 2544 16164
rect 3068 16136 3096 16204
rect 6104 16096 6132 16204
rect 1504 16068 2360 16096
rect 2700 16028 2728 16096
rect 3910 16068 4016 16096
rect 6104 16068 6684 16096
rect 8956 16068 9352 16096
rect 10060 16068 10824 16096
rect 10888 16068 11376 16096
rect 2700 16000 4200 16028
rect 4356 15892 4384 16028
rect 4632 16000 5028 16028
rect 4356 15864 5396 15892
rect 12820 15864 12940 15892
rect 1104 15728 18124 15824
rect 3528 15660 4016 15688
rect 5368 15660 6684 15688
rect 11808 15592 13032 15620
rect 4080 15524 4200 15552
rect 11808 15484 11928 15486
rect 4448 15456 4660 15484
rect 7208 15416 7236 15484
rect 7576 15456 7696 15484
rect 10336 15456 10824 15484
rect 11624 15458 12204 15484
rect 11624 15456 11836 15458
rect 11900 15456 12204 15458
rect 12544 15456 12848 15484
rect 14292 15456 15700 15484
rect 3266 15388 3372 15416
rect 4724 15388 5212 15416
rect 6932 15388 7052 15416
rect 7208 15388 7420 15416
rect 11808 15388 11854 15416
rect 7668 15320 7788 15348
rect 11624 15320 12756 15348
rect 1104 15184 18124 15280
rect 1504 15116 2084 15144
rect 3344 15116 3464 15144
rect 5736 15116 5856 15144
rect 6104 15116 7604 15144
rect 15304 15116 15608 15144
rect 1320 15048 2728 15076
rect 2332 14940 2360 15008
rect 2700 14980 2728 15048
rect 6104 15008 6132 15116
rect 10796 15048 11192 15076
rect 11716 15048 12204 15076
rect 12452 15048 13124 15076
rect 11164 15008 11192 15048
rect 3436 14980 3556 15008
rect 5920 14980 6132 15008
rect 8772 14980 9260 15008
rect 11164 14980 11836 15008
rect 12636 14994 12664 15048
rect 15120 14980 15424 15008
rect 15580 14980 15700 15008
rect 1964 14912 2084 14940
rect 2332 14912 2820 14940
rect 2792 14844 2820 14912
rect 3436 14804 3464 14980
rect 6932 14912 7052 14940
rect 8404 14912 8616 14940
rect 9232 14912 9260 14980
rect 10060 14912 10732 14940
rect 10980 14872 11008 14940
rect 12912 14872 12940 14940
rect 10980 14844 12940 14872
rect 14384 14844 14964 14872
rect 2332 14776 3464 14804
rect 7576 14776 8984 14804
rect 1104 14640 18124 14736
rect 11992 14572 12296 14600
rect 15488 14572 16436 14600
rect 12912 14504 14136 14532
rect 3344 14436 4844 14464
rect 6564 14436 6684 14464
rect 10244 14436 11100 14464
rect 11992 14436 12664 14464
rect 14108 14436 14136 14504
rect 14752 14436 16252 14464
rect 3344 14368 3372 14436
rect 8602 14368 8800 14396
rect 15856 14368 16068 14396
rect 16224 14368 16252 14436
rect 1688 14300 1808 14328
rect 2332 14300 3188 14328
rect 7208 14300 7696 14328
rect 10520 14260 10548 14328
rect 15594 14300 15700 14328
rect 1320 14232 2084 14260
rect 2148 14232 2912 14260
rect 7392 14232 9352 14260
rect 10520 14232 11468 14260
rect 15856 14232 15884 14368
rect 1104 14096 18124 14192
rect 5552 14028 6316 14056
rect 1964 13960 2912 13988
rect 15120 13960 15424 13988
rect 2056 13892 2360 13920
rect 4632 13892 4752 13920
rect 5184 13892 5764 13920
rect 5920 13892 6132 13920
rect 6840 13892 6960 13920
rect 8956 13852 8984 13920
rect 9140 13892 9352 13920
rect 11716 13892 13308 13920
rect 14660 13892 15226 13920
rect 2424 13824 2820 13852
rect 3160 13824 3740 13852
rect 7576 13824 7972 13852
rect 8956 13824 9260 13852
rect 13188 13688 13308 13716
rect 1104 13552 18124 13648
rect 11164 13484 15608 13512
rect 4540 13348 4660 13376
rect 5460 13348 6040 13376
rect 8312 13348 13860 13376
rect 5460 13308 5488 13348
rect 4172 13172 4200 13308
rect 4448 13280 5488 13308
rect 5736 13280 5856 13308
rect 4724 13212 5948 13240
rect 4724 13172 4752 13212
rect 4172 13144 4752 13172
rect 5368 13144 5764 13172
rect 5920 13144 5948 13212
rect 6012 13144 6040 13348
rect 6564 13240 6592 13308
rect 11072 13240 11100 13308
rect 11532 13280 11560 13348
rect 15028 13308 15056 13484
rect 15028 13280 15148 13308
rect 15212 13280 15424 13308
rect 15580 13280 15792 13308
rect 15396 13240 15424 13280
rect 6196 13212 6408 13240
rect 6564 13212 6960 13240
rect 9508 13212 9812 13240
rect 11072 13212 11284 13240
rect 11348 13212 12204 13240
rect 12268 13172 12296 13240
rect 15396 13212 15884 13240
rect 8588 13144 9076 13172
rect 12268 13144 12480 13172
rect 13740 13144 14228 13172
rect 1104 13008 18124 13104
rect 2424 12940 4660 12968
rect 6104 12940 6684 12968
rect 2424 12832 2452 12940
rect 1412 12804 2452 12832
rect 4356 12804 4384 12940
rect 8220 12804 8340 12832
rect 2700 12736 2820 12764
rect 4632 12736 5396 12764
rect 9140 12736 10272 12764
rect 11072 12696 11100 12764
rect 10060 12668 11100 12696
rect 13280 12696 13308 12764
rect 14476 12736 14688 12764
rect 14476 12696 14504 12736
rect 13280 12668 14504 12696
rect 4172 12600 4844 12628
rect 6472 12600 6960 12628
rect 16408 12600 16620 12628
rect 1104 12464 18124 12560
rect 3804 12396 3924 12424
rect 4632 12396 5948 12424
rect 6840 12396 7880 12424
rect 9416 12396 9720 12424
rect 10612 12288 10640 12424
rect 1780 12260 2176 12288
rect 2792 12260 2912 12288
rect 9968 12260 10640 12288
rect 12360 12260 14504 12288
rect 14752 12260 14964 12288
rect 1688 12152 1716 12220
rect 2148 12192 2176 12260
rect 2746 12192 4016 12220
rect 7944 12192 9352 12220
rect 9968 12192 9996 12260
rect 12452 12192 12848 12220
rect 12912 12192 13400 12220
rect 1688 12124 2268 12152
rect 2746 12084 2774 12192
rect 12452 12152 12480 12192
rect 12912 12152 12940 12192
rect 13740 12152 13768 12220
rect 13924 12192 14228 12220
rect 4632 12124 4752 12152
rect 5828 12124 7328 12152
rect 12360 12124 12480 12152
rect 12544 12124 12940 12152
rect 13004 12124 13584 12152
rect 13740 12124 14780 12152
rect 2056 12056 2774 12084
rect 11348 12056 12756 12084
rect 1104 11920 18124 12016
rect 4632 11852 4844 11880
rect 4908 11852 5488 11880
rect 5736 11852 5856 11880
rect 11532 11852 12112 11880
rect 16960 11812 16988 11880
rect 17144 11852 17540 11880
rect 17144 11812 17172 11852
rect 4724 11784 5304 11812
rect 14490 11784 15056 11812
rect 16960 11784 17172 11812
rect 17236 11784 17724 11812
rect 2976 11716 3556 11744
rect 4816 11716 5120 11744
rect 5368 11716 7972 11744
rect 15120 11716 15792 11744
rect 16960 11716 17540 11744
rect 5368 11676 5396 11716
rect 16960 11676 16988 11716
rect 3988 11648 5396 11676
rect 4080 11580 4568 11608
rect 13004 11540 13032 11676
rect 13280 11648 13400 11676
rect 13648 11648 14596 11676
rect 16592 11648 16988 11676
rect 14568 11540 14596 11648
rect 14844 11580 16712 11608
rect 5184 11512 5304 11540
rect 13004 11512 14504 11540
rect 14568 11512 17080 11540
rect 1104 11376 18124 11472
rect 4724 11308 6776 11336
rect 8404 11308 8616 11336
rect 16224 11240 16712 11268
rect 16684 11200 16712 11240
rect 1412 11172 3832 11200
rect 5920 11172 6868 11200
rect 7116 11172 9536 11200
rect 9692 11172 14504 11200
rect 14752 11172 14872 11200
rect 16684 11172 17356 11200
rect 9232 11104 9352 11132
rect 12084 11104 12388 11132
rect 12544 11064 12572 11132
rect 1688 11036 1808 11064
rect 9048 11036 9260 11064
rect 12176 11036 12572 11064
rect 16868 11036 17356 11064
rect 9232 10968 9260 11036
rect 11440 10968 12020 10996
rect 1104 10832 18124 10928
rect 1504 10764 2084 10792
rect 2148 10764 2268 10792
rect 2332 10764 2820 10792
rect 3436 10764 8800 10792
rect 10704 10764 10824 10792
rect 11808 10764 13308 10792
rect 13372 10764 13676 10792
rect 1964 10656 1992 10724
rect 2332 10696 2360 10764
rect 4816 10696 4936 10724
rect 8772 10696 8800 10764
rect 12912 10696 13216 10724
rect 1964 10628 2452 10656
rect 3358 10628 3556 10656
rect 5184 10628 5396 10656
rect 5552 10628 5856 10656
rect 10704 10628 10824 10656
rect 13004 10628 13584 10656
rect 3160 10560 3280 10588
rect 4540 10560 5488 10588
rect 6196 10560 6684 10588
rect 6748 10560 11560 10588
rect 12084 10560 12480 10588
rect 14936 10560 16712 10588
rect 8128 10492 8340 10520
rect 10980 10492 13032 10520
rect 1104 10288 18124 10384
rect 8680 10220 8984 10248
rect 4816 10084 5580 10112
rect 5644 10084 5948 10112
rect 8312 10084 8524 10112
rect 11992 10084 12848 10112
rect 1964 10016 3832 10044
rect 5460 10016 5764 10044
rect 5920 10016 5948 10084
rect 8496 10016 8524 10084
rect 9600 10016 10732 10044
rect 12544 10016 12664 10044
rect 12820 10016 12848 10084
rect 17328 10084 17632 10112
rect 17328 10044 17356 10084
rect 14476 10016 14688 10044
rect 16684 10016 17356 10044
rect 3896 9880 4200 9908
rect 16408 9880 16528 9908
rect 1104 9744 18124 9840
rect 4632 9676 4752 9704
rect 16684 9676 16896 9704
rect 16960 9636 16988 9704
rect 2792 9608 3188 9636
rect 6840 9568 6868 9636
rect 8220 9608 9168 9636
rect 1872 9540 1992 9568
rect 6656 9540 6868 9568
rect 7760 9540 7972 9568
rect 8220 9540 8248 9608
rect 8588 9500 8616 9568
rect 9140 9540 9168 9608
rect 9876 9608 10732 9636
rect 11716 9608 11928 9636
rect 16776 9608 17172 9636
rect 9876 9568 9904 9608
rect 10704 9568 10732 9608
rect 9232 9540 9904 9568
rect 10520 9540 10640 9568
rect 10704 9540 12112 9568
rect 15396 9540 15516 9568
rect 17052 9540 17540 9568
rect 9232 9500 9260 9540
rect 2884 9364 2912 9500
rect 6380 9472 6868 9500
rect 8312 9472 8524 9500
rect 8588 9472 9260 9500
rect 8588 9432 8616 9472
rect 7024 9404 8616 9432
rect 14752 9404 17264 9432
rect 2884 9336 4568 9364
rect 7852 9336 8524 9364
rect 10060 9336 10364 9364
rect 1104 9200 18124 9296
rect 4080 9132 5672 9160
rect 10796 9132 13216 9160
rect 4080 9024 4108 9132
rect 2056 8996 4108 9024
rect 1320 8928 1808 8956
rect 2056 8928 2084 8996
rect 2700 8888 2728 8956
rect 2884 8928 3004 8956
rect 4080 8928 4108 8996
rect 8956 8996 11468 9024
rect 8956 8956 8984 8996
rect 4264 8888 4292 8956
rect 8588 8928 8984 8956
rect 2700 8860 3280 8888
rect 4264 8860 4752 8888
rect 2056 8792 2544 8820
rect 4724 8792 4752 8860
rect 4908 8820 4936 8888
rect 12558 8860 13124 8888
rect 13188 8820 13216 9132
rect 16224 8956 16252 9024
rect 16132 8928 16528 8956
rect 4908 8792 5764 8820
rect 13188 8792 15424 8820
rect 1104 8656 18124 8752
rect 1320 8588 1808 8616
rect 1872 8588 2268 8616
rect 7852 8588 8340 8616
rect 8404 8588 9536 8616
rect 8404 8548 8432 8588
rect 9600 8548 9628 8616
rect 10612 8588 12848 8616
rect 16408 8588 16712 8616
rect 2148 8480 2176 8548
rect 4632 8520 4936 8548
rect 5920 8520 7236 8548
rect 7760 8520 8432 8548
rect 9140 8520 9628 8548
rect 9784 8520 10088 8548
rect 5920 8480 5948 8520
rect 1688 8452 2176 8480
rect 3082 8452 3280 8480
rect 3896 8452 4016 8480
rect 4448 8452 5948 8480
rect 6104 8412 6132 8480
rect 6380 8452 6500 8480
rect 8864 8452 9996 8480
rect 10888 8466 10916 8588
rect 11440 8520 14504 8548
rect 11532 8452 11652 8480
rect 16224 8452 16528 8480
rect 4816 8384 5396 8412
rect 6104 8384 7052 8412
rect 10704 8384 10824 8412
rect 15672 8384 16712 8412
rect 1504 8316 1716 8344
rect 1104 8112 18124 8208
rect 2976 8044 3188 8072
rect 3252 8044 3924 8072
rect 4632 7908 5672 7936
rect 14476 7908 15976 7936
rect 6288 7840 6500 7868
rect 12728 7800 12756 7868
rect 12912 7840 13308 7868
rect 16776 7840 17080 7868
rect 17328 7840 17632 7868
rect 5644 7772 6132 7800
rect 12728 7772 13032 7800
rect 14384 7772 14490 7800
rect 4724 7704 6040 7732
rect 6104 7704 6132 7772
rect 12176 7704 12296 7732
rect 14200 7704 14320 7732
rect 1104 7568 18124 7664
rect 4540 7500 4660 7528
rect 7024 7460 7052 7528
rect 8680 7500 9812 7528
rect 5736 7432 6776 7460
rect 7024 7432 7788 7460
rect 1964 7364 2084 7392
rect 7760 7364 7788 7432
rect 8036 7432 8616 7460
rect 9522 7432 10088 7460
rect 8036 7364 8064 7432
rect 9876 7364 10180 7392
rect 10980 7364 11284 7392
rect 11440 7364 11560 7392
rect 14292 7364 15424 7392
rect 1104 7024 18124 7120
rect 6472 6956 6665 6984
rect 4080 6888 4660 6916
rect 11072 6888 11836 6916
rect 4080 6848 4108 6888
rect 1412 6820 4108 6848
rect 4816 6820 4936 6848
rect 5736 6820 6132 6848
rect 6288 6820 7052 6848
rect 8128 6820 9260 6848
rect 3988 6752 5580 6780
rect 5644 6712 5672 6780
rect 3266 6684 3924 6712
rect 4264 6684 5304 6712
rect 5552 6684 5672 6712
rect 4632 6616 4752 6644
rect 5552 6616 5580 6684
rect 5736 6644 5764 6820
rect 6104 6752 6132 6820
rect 9232 6752 9260 6820
rect 11256 6820 12296 6848
rect 10336 6644 10364 6780
rect 11256 6752 11284 6820
rect 11624 6752 12572 6780
rect 14292 6752 14412 6780
rect 5644 6616 5764 6644
rect 8588 6616 9076 6644
rect 10336 6616 11376 6644
rect 11440 6616 13676 6644
rect 1104 6480 18124 6576
rect 2056 6412 2728 6440
rect 5552 6412 6960 6440
rect 8128 6412 8248 6440
rect 8404 6412 11192 6440
rect 3988 6344 4200 6372
rect 5644 6344 5948 6372
rect 3988 6276 4016 6344
rect 6932 6304 6960 6412
rect 8404 6372 8432 6412
rect 7760 6344 8432 6372
rect 10428 6344 11468 6372
rect 6932 6276 7604 6304
rect 7944 6276 8248 6304
rect 8312 6276 8360 6304
rect 10336 6276 10640 6304
rect 10704 6276 10824 6304
rect 11900 6276 11965 6304
rect 12084 6276 12388 6304
rect 10612 6236 10640 6276
rect 11900 6236 11928 6276
rect 5552 6208 5856 6236
rect 10612 6208 10916 6236
rect 11348 6208 12848 6236
rect 5460 6140 7420 6168
rect 10060 6140 10272 6168
rect 5736 6072 5856 6100
rect 12452 6072 12664 6100
rect 14568 6072 15056 6100
rect 1104 5936 18124 6032
rect 4080 5800 7052 5828
rect 13096 5800 13308 5828
rect 4080 5760 4108 5800
rect 1596 5732 4108 5760
rect 1596 5692 1624 5732
rect 1412 5664 1624 5692
rect 1872 5596 1992 5624
rect 3252 5596 3832 5624
rect 3252 5556 3280 5596
rect 4816 5556 4844 5692
rect 5276 5664 5304 5800
rect 10060 5732 10548 5760
rect 10796 5732 11376 5760
rect 10796 5664 10824 5732
rect 13464 5664 14228 5692
rect 14292 5664 14582 5692
rect 11256 5556 11284 5624
rect 13464 5596 13492 5664
rect 2148 5528 3280 5556
rect 3344 5528 4844 5556
rect 8496 5528 8708 5556
rect 9048 5528 10548 5556
rect 11256 5528 12296 5556
rect 13004 5528 13124 5556
rect 1104 5392 18124 5488
rect 1504 5324 2268 5352
rect 2700 5324 2912 5352
rect 3436 5324 4752 5352
rect 5368 5324 6132 5352
rect 13832 5324 14504 5352
rect 1504 5216 1532 5324
rect 2516 5256 3280 5284
rect 1320 5188 1532 5216
rect 1780 5148 1808 5216
rect 2056 5188 3004 5216
rect 3436 5188 3464 5324
rect 4356 5256 4660 5284
rect 5842 5256 6224 5284
rect 6840 5256 8248 5284
rect 11348 5256 11468 5284
rect 4356 5188 4384 5256
rect 6104 5188 6578 5216
rect 7760 5188 7880 5216
rect 8220 5188 8248 5256
rect 9968 5202 10442 5216
rect 9968 5188 10456 5202
rect 14292 5188 14688 5216
rect 14844 5188 15056 5216
rect 6104 5148 6132 5188
rect 1780 5120 2360 5148
rect 5644 5120 6132 5148
rect 6656 5080 6684 5148
rect 9968 5120 9996 5188
rect 5828 5052 6684 5080
rect 10428 5080 10456 5188
rect 10520 5120 10916 5148
rect 10428 5052 10640 5080
rect 1104 4848 18124 4944
rect 5368 4780 5580 4808
rect 9232 4780 9352 4808
rect 9508 4780 9904 4808
rect 10704 4780 10916 4808
rect 4172 4712 4660 4740
rect 4816 4712 6500 4740
rect 4172 4644 4200 4712
rect 5736 4644 5856 4672
rect 10520 4644 10916 4672
rect 5552 4576 5672 4604
rect 6288 4468 6316 4604
rect 8220 4576 9996 4604
rect 10612 4576 10732 4604
rect 11440 4576 11928 4604
rect 13648 4576 14136 4604
rect 7852 4508 7972 4536
rect 8220 4468 8248 4576
rect 13924 4508 14412 4536
rect 6288 4440 8248 4468
rect 15764 4440 15884 4468
rect 1104 4304 18124 4400
rect 2746 4236 5396 4264
rect 6380 4236 6868 4264
rect 6932 4236 7788 4264
rect 2746 4196 2774 4236
rect 6932 4196 6960 4236
rect 1780 4168 2774 4196
rect 4816 4168 5488 4196
rect 6656 4168 6960 4196
rect 7116 4168 7604 4196
rect 6656 4128 6684 4168
rect 4586 4100 4936 4128
rect 5184 4100 6684 4128
rect 6748 4100 7420 4128
rect 7668 4100 7774 4128
rect 9600 4100 11008 4128
rect 13004 4060 13032 4128
rect 13188 4100 13768 4128
rect 14384 4100 14872 4128
rect 14936 4100 15424 4128
rect 2148 4032 2360 4060
rect 12820 4032 13584 4060
rect 2148 3896 2176 4032
rect 4080 3964 4292 3992
rect 4816 3964 5028 3992
rect 6472 3964 6592 3992
rect 2332 3896 2728 3924
rect 10612 3896 10916 3924
rect 1104 3760 18124 3856
rect 7944 3692 8248 3720
rect 9968 3692 10548 3720
rect 9140 3624 10272 3652
rect 1688 3556 2176 3584
rect 4264 3556 4660 3584
rect 5000 3556 5856 3584
rect 9140 3516 9168 3624
rect 10520 3584 10548 3692
rect 2976 3488 3556 3516
rect 3804 3502 4554 3516
rect 3804 3488 4568 3502
rect 4540 3448 4568 3488
rect 5644 3448 5672 3516
rect 8956 3488 9168 3516
rect 9232 3556 10364 3584
rect 10520 3556 10640 3584
rect 11532 3556 11928 3584
rect 9232 3488 9260 3556
rect 2898 3420 3464 3448
rect 4540 3420 5672 3448
rect 9324 3420 9720 3448
rect 9968 3420 10180 3448
rect 10336 3380 10364 3556
rect 11532 3502 11560 3556
rect 13740 3488 14412 3516
rect 14844 3488 14964 3516
rect 14384 3448 14412 3488
rect 10520 3420 11928 3448
rect 13832 3420 14320 3448
rect 14384 3420 14504 3448
rect 14660 3420 15976 3448
rect 1964 3352 3188 3380
rect 8680 3352 9536 3380
rect 9784 3352 10088 3380
rect 10336 3352 13768 3380
rect 13924 3352 14228 3380
rect 14476 3352 14504 3420
rect 14844 3352 14964 3380
rect 1104 3216 18124 3312
rect 2056 3148 6224 3176
rect 9508 3148 13676 3176
rect 2056 3040 2084 3148
rect 4080 3108 4108 3148
rect 1412 3012 2084 3040
rect 3988 3080 4108 3108
rect 4172 3080 4292 3108
rect 5474 3080 6040 3108
rect 7484 3080 7880 3108
rect 3988 3012 4016 3080
rect 9508 3040 9536 3148
rect 12268 3080 13400 3108
rect 13556 3080 13860 3108
rect 13556 3040 13584 3080
rect 6104 3012 6316 3040
rect 9416 3012 9536 3040
rect 11256 3012 11652 3040
rect 13280 3012 13584 3040
rect 6288 2972 6316 3012
rect 6288 2944 7236 2972
rect 11256 2944 11284 3012
rect 15396 2944 15608 2972
rect 1104 2672 18124 2768
rect 2424 2604 2544 2632
rect 7116 2604 7328 2632
rect 7576 2604 7696 2632
rect 12360 2604 13032 2632
rect 12452 2536 14412 2564
rect 8036 2468 8248 2496
rect 9048 2468 9168 2496
rect 2516 2400 2636 2428
rect 7668 2400 7880 2428
rect 12452 2400 12480 2536
rect 12820 2468 12940 2496
rect 13004 2468 13768 2496
rect 14292 2468 14688 2496
rect 13004 2428 13032 2468
rect 12728 2400 13032 2428
rect 13096 2400 14872 2428
rect 15594 2400 15792 2428
rect 1104 2128 18124 2224
<< metal2 >>
rect 1504 16068 1532 19802
rect 1964 18244 1992 18680
rect 1596 17564 1624 18068
rect 1688 16136 1716 16504
rect 1780 15524 1808 17728
rect 2240 17292 2268 19122
rect 2792 17836 2820 20482
rect 2976 17564 3004 18204
rect 3160 17836 3188 18068
rect 3344 17224 3372 18204
rect 2148 16204 2176 16504
rect 2884 16266 2912 16640
rect 2792 16238 2912 16266
rect 2792 16204 2820 16238
rect 2056 15116 2084 15416
rect 1320 14232 1348 15076
rect 1688 13348 1716 14328
rect 1964 13960 1992 14940
rect 1412 11172 1440 13308
rect 1504 10764 1532 12220
rect 1780 10696 1808 11064
rect 1964 10696 1992 12220
rect 2056 10554 2084 13920
rect 2148 11036 2176 11540
rect 1964 10526 2084 10554
rect 1872 9132 1900 9568
rect 1320 8588 1348 8956
rect 1688 7908 1716 8344
rect 1412 6820 1440 7868
rect 1320 4134 1348 5216
rect 1412 3012 1440 5692
rect 1872 5256 1900 6304
rect 1964 5794 1992 10526
rect 2056 8520 2084 8820
rect 2148 8520 2176 9500
rect 2240 8588 2268 14260
rect 2332 13892 2360 16096
rect 2884 15694 2912 16238
rect 2976 15586 3004 17184
rect 3252 16068 3280 16436
rect 2884 15558 3004 15586
rect 2884 14232 2912 15558
rect 3344 15116 3372 15416
rect 3344 13892 3372 14396
rect 2792 13280 2820 13852
rect 3160 13484 3188 13852
rect 2792 12260 2820 12764
rect 2792 10764 2820 11540
rect 3160 10560 3188 11676
rect 3436 10764 3464 21162
rect 3620 17224 3648 18340
rect 3804 16680 3832 18680
rect 4632 17224 4660 18612
rect 4540 16612 4660 16640
rect 3988 15660 4016 16572
rect 4172 16204 4200 16436
rect 4540 16374 4568 16612
rect 4724 16574 4752 18680
rect 4816 17632 4844 18748
rect 5460 16612 5488 18408
rect 5552 16680 5580 18340
rect 5644 17564 5672 18136
rect 5736 17490 5764 18272
rect 5644 17462 5764 17490
rect 5644 16612 5672 17462
rect 4724 16546 4844 16574
rect 4080 15524 4108 16028
rect 4632 15456 4660 16504
rect 3528 13824 3556 14396
rect 4172 13818 4200 14362
rect 4080 13790 4200 13818
rect 4080 13410 4108 13790
rect 4080 13382 4200 13410
rect 4172 13280 4200 13382
rect 4632 13348 4660 13920
rect 3804 12396 3832 12832
rect 4632 12396 4660 13240
rect 2976 8044 3004 8956
rect 3252 8044 3280 8888
rect 2148 7500 2176 7800
rect 3528 6956 3556 11744
rect 3988 11648 4016 12220
rect 4080 11172 4108 11608
rect 4172 9608 4200 9908
rect 4632 9574 4660 11880
rect 4724 11308 4752 15416
rect 4816 12600 4844 16546
rect 6012 16204 6040 17184
rect 6104 17156 6132 17524
rect 6196 16204 6224 18272
rect 6472 17632 6500 18068
rect 5000 15524 5028 16028
rect 5368 15660 5396 15892
rect 5736 15116 5764 16096
rect 5828 13960 5856 14328
rect 5368 12736 5396 13172
rect 4816 10696 4844 11744
rect 5184 11104 5212 11540
rect 5276 11098 5304 11812
rect 5460 11098 5488 13376
rect 5736 13002 5764 13920
rect 5736 12974 5856 13002
rect 5736 11852 5764 12832
rect 5828 12124 5856 12974
rect 5920 11172 5948 12424
rect 6104 11716 6132 15008
rect 6656 14436 6684 17728
rect 6748 16068 6776 17524
rect 7024 16612 7052 17116
rect 7116 16544 7144 16980
rect 7484 16574 7512 18748
rect 8220 18312 8248 18612
rect 7760 17660 7788 18068
rect 8772 17768 8800 18204
rect 7668 17632 7788 17660
rect 7668 17088 7696 17632
rect 8496 17292 8524 17660
rect 6288 14028 6316 14328
rect 6932 13892 6960 15416
rect 7024 14504 7052 14940
rect 7208 13892 7236 14328
rect 7300 13382 7328 15484
rect 7392 14232 7420 16572
rect 7484 16546 7604 16574
rect 7576 15116 7604 16546
rect 7760 16544 7788 17252
rect 8772 16574 8800 17592
rect 9232 17054 9260 17524
rect 9324 17156 9352 17524
rect 8772 16546 8892 16574
rect 8864 16000 8892 16546
rect 9324 16068 9352 16980
rect 9416 16612 9444 18204
rect 9508 17292 9536 17592
rect 9692 17224 9720 18204
rect 9416 16204 9444 16504
rect 10060 16068 10088 18748
rect 10428 18312 10456 18612
rect 10612 17728 10640 17762
rect 10612 17700 10824 17728
rect 11164 17700 11192 18068
rect 10520 17224 10548 17524
rect 10612 17292 10640 17700
rect 10704 16748 10732 17592
rect 10796 17156 10824 17700
rect 11348 17224 11376 17660
rect 10152 16204 10180 16504
rect 7668 15048 7696 15348
rect 10244 15048 10272 15348
rect 10796 15048 10824 16572
rect 7576 14368 7604 14804
rect 8496 14436 8524 14940
rect 8772 14368 8800 15008
rect 6656 12730 6684 13308
rect 6656 12702 6776 12730
rect 6748 12260 6776 12702
rect 6840 12396 6868 12832
rect 6932 12192 6960 13240
rect 7944 12872 7972 13852
rect 8312 12804 8340 13376
rect 8588 12872 8616 13172
rect 9140 12736 9168 14464
rect 10060 14436 10088 14940
rect 11072 14436 11100 14872
rect 11348 14844 11376 17116
rect 9232 13960 9260 14396
rect 11256 14300 11284 14804
rect 9232 12838 9260 13852
rect 9324 12628 9352 14260
rect 11440 14232 11468 15416
rect 11164 13280 11192 13512
rect 11256 13246 11376 13274
rect 9140 12600 9352 12628
rect 5276 11070 5396 11098
rect 5460 11070 5672 11098
rect 4724 9676 4752 10656
rect 5368 9948 5396 11070
rect 5552 10588 5580 10996
rect 5460 10560 5580 10588
rect 5552 10084 5580 10560
rect 5460 9574 5488 10044
rect 4540 9438 4660 9466
rect 4540 9336 4568 9438
rect 3896 8452 3924 8888
rect 2056 6412 2084 6712
rect 4172 6344 4200 6916
rect 4264 6344 4292 6712
rect 1964 5766 2084 5794
rect 1964 5256 1992 5624
rect 1688 2774 1716 4196
rect 1780 4168 1808 5216
rect 2056 5188 2084 5766
rect 2148 5256 2176 6236
rect 2332 5120 2360 5352
rect 2884 5324 2912 5624
rect 1964 2400 1992 4128
rect 2148 3556 2176 3924
rect 2332 3080 2360 3924
rect 2148 2400 2176 2802
rect 2516 2604 2544 4128
rect 2608 2400 2636 4196
rect 2976 3488 3004 5216
rect 3620 5188 3648 5556
rect 4632 5256 4660 9438
rect 4724 7704 4752 8820
rect 4816 6820 4844 7800
rect 5368 7772 5396 8412
rect 5644 7772 5672 11070
rect 5828 10220 5856 10656
rect 6380 10628 6408 11200
rect 5736 7976 5764 8820
rect 6012 8588 6040 8956
rect 5920 7840 5948 8480
rect 6380 8452 6408 9500
rect 6472 7840 6500 9364
rect 4724 6344 4752 6644
rect 5460 6140 5488 6712
rect 5552 6412 5580 6780
rect 5644 6344 5672 6780
rect 4632 4712 4660 5148
rect 4724 5114 4752 5692
rect 4724 5086 4844 5114
rect 4816 4712 4844 5086
rect 4632 4128 4660 4604
rect 4448 4100 4660 4128
rect 3436 2604 3464 3040
rect 3528 2400 3556 3516
rect 3804 2944 3832 3516
rect 4080 3108 4108 3992
rect 4632 3556 4660 4100
rect 4816 3964 4844 4604
rect 4908 3454 4936 4128
rect 5368 4100 5396 5352
rect 5552 4780 5580 6236
rect 5736 5664 5764 7460
rect 5828 6208 5856 6780
rect 5644 4576 5672 5148
rect 5828 4644 5856 6100
rect 5920 5086 5948 6780
rect 6104 5324 6132 7732
rect 6748 7432 6776 11336
rect 6840 8452 6868 9636
rect 7024 7562 7052 11744
rect 7944 11716 7972 12220
rect 7852 11036 7880 11540
rect 7116 10220 7144 10724
rect 8312 10084 8340 11744
rect 8404 10016 8432 11676
rect 8956 10220 8984 11064
rect 9048 10146 9076 11064
rect 8956 10118 9076 10146
rect 7760 7806 7788 9568
rect 8956 9540 8984 10118
rect 7852 8860 7880 9364
rect 8312 8588 8340 8888
rect 8496 8452 8524 9500
rect 6932 7534 7052 7562
rect 6472 6956 6500 7324
rect 6196 4780 6224 5284
rect 5460 3692 5488 4196
rect 4080 3080 4200 3108
rect 5736 2944 5764 3584
rect 6196 3148 6224 3516
rect 6288 3012 6316 6440
rect 6380 5800 6408 6780
rect 6932 6412 6960 7534
rect 7024 7500 7052 7534
rect 7024 6820 7052 7392
rect 6840 5256 6868 5828
rect 7392 5120 7420 7392
rect 7668 6684 7696 7188
rect 7484 4508 7512 6100
rect 7668 5188 7696 5250
rect 6380 2366 6408 4264
rect 7760 4236 7788 6372
rect 7944 5732 7972 7800
rect 8312 6474 8340 7324
rect 8404 6820 8432 7868
rect 8588 7432 8616 8956
rect 9140 8520 9168 12600
rect 9692 12396 9720 12832
rect 9784 12396 9812 13240
rect 11256 13212 11284 13246
rect 10060 12192 10088 12696
rect 10612 12396 10640 12832
rect 11348 12056 11376 13246
rect 11532 12434 11560 16096
rect 11624 15320 11652 18306
rect 11808 17224 11836 17524
rect 11992 17292 12020 17524
rect 11808 15388 11836 16980
rect 12544 16748 12572 17252
rect 11808 13892 11836 15008
rect 11992 14572 12020 15416
rect 12176 15048 12204 15484
rect 12452 14368 12480 15076
rect 12544 14436 12572 14940
rect 12728 14368 12756 15348
rect 12820 14572 12848 15484
rect 12912 14504 12940 15892
rect 11440 12406 11560 12434
rect 9232 10084 9260 11676
rect 9968 10084 9996 11064
rect 10704 10764 10732 11064
rect 9324 9608 9352 10044
rect 9600 8996 9628 10044
rect 9232 8384 9260 8888
rect 8680 7500 8708 7868
rect 9324 6752 9352 7528
rect 9876 7364 9904 9568
rect 9968 8860 9996 9364
rect 10060 8520 10088 9364
rect 10612 8588 10640 9568
rect 10704 8384 10732 9500
rect 10796 9132 10824 10656
rect 11440 10588 11468 12406
rect 11624 12124 11652 13852
rect 12084 11852 12112 12152
rect 12176 11716 12204 13240
rect 12452 12328 12480 13172
rect 11808 10662 11836 11132
rect 12360 11104 12388 12152
rect 12544 11716 12572 12152
rect 12820 12056 12848 13512
rect 13004 13484 13032 15620
rect 13096 15048 13124 16980
rect 14292 15456 14320 16640
rect 13188 15048 13216 15348
rect 14200 15048 14228 15348
rect 14384 14436 14412 14872
rect 14660 14464 14688 14804
rect 14660 14436 14780 14464
rect 14660 13892 14688 14436
rect 13280 13212 13308 13716
rect 13372 12192 13400 12764
rect 13832 12668 13860 13376
rect 15212 13280 15240 15144
rect 14108 12124 14136 12832
rect 14200 12192 14228 13172
rect 11440 10560 11560 10588
rect 10980 10084 11008 10520
rect 11348 7500 11376 8888
rect 10336 6752 10364 6882
rect 10704 6820 10732 7392
rect 8220 6446 8340 6474
rect 8220 6412 8248 6446
rect 8588 6344 8616 6644
rect 10612 6412 10640 6780
rect 11256 6752 11284 7392
rect 11440 7364 11468 9024
rect 11348 6616 11468 6644
rect 11164 6338 11192 6440
rect 11348 6338 11376 6616
rect 11164 6310 11376 6338
rect 8036 5188 8064 5692
rect 8312 5222 8340 6304
rect 10336 6174 10364 6304
rect 10060 5732 10088 6168
rect 8496 5256 8524 5556
rect 8220 4644 8248 5216
rect 9232 4780 9260 5284
rect 9508 4780 9536 5624
rect 10520 5120 10548 5556
rect 6472 3556 6500 3992
rect 6656 2400 6684 4128
rect 6748 2468 6776 3040
rect 6932 3012 6960 4128
rect 7116 2604 7144 3448
rect 7208 2400 7236 2972
rect 7576 2604 7604 4196
rect 7668 2400 7696 4128
rect 7852 3080 7880 4536
rect 8220 2468 8248 4060
rect 8680 3080 8708 3380
rect 8956 1414 8984 3516
rect 9600 3488 9628 4604
rect 10612 4576 10640 5080
rect 10704 4780 10732 6304
rect 9140 2468 9168 2972
rect 9692 2400 9720 3448
rect 9784 3080 9812 3380
rect 9968 2400 9996 3720
rect 10244 3352 10272 3652
rect 10612 3108 10640 3924
rect 10796 3148 10824 5692
rect 10888 5664 10916 6236
rect 11164 5664 11192 6310
rect 11348 5732 11376 6236
rect 10888 4644 10916 5148
rect 11440 4576 11468 6372
rect 11532 5256 11560 10560
rect 11992 10084 12020 10996
rect 12912 10696 12940 11132
rect 13372 11104 13400 11676
rect 12452 10146 12480 10588
rect 13004 10220 13032 10656
rect 12452 10118 12572 10146
rect 12544 10016 12572 10118
rect 11716 9608 11744 9976
rect 11808 6888 11836 7324
rect 12084 6276 12112 9568
rect 12820 8588 12848 8820
rect 12268 7432 12296 7732
rect 12544 6752 12572 7732
rect 11624 4644 11652 5624
rect 12636 5596 12664 6100
rect 12268 4576 12296 5556
rect 12820 5324 12848 6236
rect 13004 5528 13032 7800
rect 13280 6752 13308 7868
rect 13096 5800 13124 6236
rect 13280 4168 13308 4604
rect 13464 4576 13492 5624
rect 13648 5556 13676 11676
rect 14476 11172 14504 12764
rect 14936 12260 14964 12764
rect 15304 12192 15332 13444
rect 15396 12260 15424 15008
rect 15488 14572 15516 15008
rect 15580 13484 15608 15144
rect 15672 15008 15700 15484
rect 15672 14980 15792 15008
rect 15672 14300 15700 14804
rect 15672 12872 15700 13172
rect 14752 11852 14780 12152
rect 14844 11172 14872 11608
rect 14936 10084 14964 10588
rect 14476 7908 14504 10044
rect 14752 8996 14780 9432
rect 14200 6276 14228 6644
rect 10520 3080 10640 3108
rect 11624 3012 11652 3516
rect 11716 3012 11744 3584
rect 11900 3080 11928 3448
rect 12360 2604 12388 3448
rect 12452 734 12480 2428
rect 12820 54 12848 4060
rect 13556 4032 13584 5556
rect 13648 5528 13768 5556
rect 13372 3080 13400 3448
rect 12912 2468 12940 3040
rect 13648 3012 13676 4604
rect 13740 2468 13768 5528
rect 13832 5324 13860 5624
rect 14292 5188 14320 7732
rect 14384 7500 14412 7800
rect 14384 4100 14412 7392
rect 15396 7364 15424 11744
rect 15764 11716 15792 14980
rect 15856 13892 15884 14260
rect 15488 10764 15516 11064
rect 15856 10526 15884 13240
rect 16592 11104 16620 12628
rect 16868 11036 16896 11744
rect 17052 11512 17080 11880
rect 17328 11172 17356 11676
rect 17328 10560 17356 11064
rect 17420 10220 17448 10656
rect 15580 9608 15608 9976
rect 16500 9466 16528 9908
rect 16684 9676 16712 10044
rect 17512 10016 17540 11880
rect 16500 9438 16620 9466
rect 15488 8588 15516 8888
rect 16132 8452 16160 8956
rect 16592 8922 16620 9438
rect 16500 8894 16620 8922
rect 16500 8452 16528 8894
rect 16684 8588 16712 9568
rect 15672 7772 15700 8412
rect 16776 7840 16804 9636
rect 17144 9574 17172 9636
rect 17420 7908 17448 8480
rect 17512 8384 17540 9568
rect 17604 7840 17632 11642
rect 15028 5188 15056 6100
rect 13832 3080 13860 3448
rect 13924 3080 13952 3380
rect 14292 2468 14320 3448
rect 14384 2536 14412 3380
rect 14844 2400 14872 4128
rect 15396 4100 15424 4536
rect 14936 3080 14964 3380
rect 15488 2468 15516 2972
rect 15764 2400 15792 4468
rect 15948 3148 15976 3448
<< metal3 >>
rect 0 21178 800 21208
rect 0 21118 3480 21178
rect 0 21088 800 21118
rect 0 20498 800 20528
rect 0 20438 2836 20498
rect 0 20408 800 20438
rect 0 19818 800 19848
rect 0 19758 1548 19818
rect 0 19728 800 19758
rect 0 19138 800 19168
rect 0 19078 2284 19138
rect 0 19048 800 19078
rect 4170 19007 4566 19073
rect 10170 19007 10566 19073
rect 16170 19007 16566 19073
rect 0 18458 800 18488
rect 4910 18463 5306 18529
rect 10910 18463 11306 18529
rect 16910 18463 17306 18529
rect 0 18398 3434 18458
rect 0 18368 800 18398
rect 3374 18322 3434 18398
rect 3374 18262 11668 18322
rect 4170 17919 4566 17985
rect 10170 17919 10566 17985
rect 16170 17919 16566 17985
rect 0 17778 800 17808
rect 0 17718 10656 17778
rect 0 17688 800 17718
rect 4910 17375 5306 17441
rect 10910 17375 11306 17441
rect 16910 17375 17306 17441
rect 0 17098 800 17128
rect 0 17038 9276 17098
rect 0 17008 800 17038
rect 4170 16831 4566 16897
rect 10170 16831 10566 16897
rect 16170 16831 16566 16897
rect 0 16418 800 16448
rect 0 16358 4584 16418
rect 0 16328 800 16358
rect 4910 16287 5306 16353
rect 10910 16287 11306 16353
rect 16910 16287 17306 16353
rect 0 15738 800 15768
rect 4170 15743 4566 15809
rect 10170 15743 10566 15809
rect 16170 15743 16566 15809
rect 0 15678 2928 15738
rect 0 15648 800 15678
rect 4910 15199 5306 15265
rect 10910 15199 11306 15265
rect 16910 15199 17306 15265
rect 0 15058 800 15088
rect 0 14998 1364 15058
rect 0 14968 800 14998
rect 4170 14655 4566 14721
rect 10170 14655 10566 14721
rect 16170 14655 16566 14721
rect 0 14378 800 14408
rect 0 14318 4216 14378
rect 0 14288 800 14318
rect 4910 14111 5306 14177
rect 10910 14111 11306 14177
rect 16910 14111 17306 14177
rect 0 13698 800 13728
rect 0 13638 3434 13698
rect 0 13608 800 13638
rect 3374 13426 3434 13638
rect 4170 13567 4566 13633
rect 10170 13567 10566 13633
rect 16170 13567 16566 13633
rect 3374 13366 7344 13426
rect 0 13018 800 13048
rect 4910 13023 5306 13089
rect 10910 13023 11306 13089
rect 16910 13023 17306 13089
rect 0 12958 3066 13018
rect 0 12928 800 12958
rect 3006 12882 3066 12958
rect 3006 12822 9276 12882
rect 4170 12479 4566 12545
rect 10170 12479 10566 12545
rect 16170 12479 16566 12545
rect 0 12338 800 12368
rect 0 12278 11392 12338
rect 0 12248 800 12278
rect 4910 11935 5306 12001
rect 10910 11935 11306 12001
rect 16910 11935 17306 12001
rect 0 11658 800 11688
rect 18507 11658 19307 11688
rect 0 11598 1548 11658
rect 17036 11598 19307 11658
rect 0 11568 800 11598
rect 18507 11568 19307 11598
rect 4170 11391 4566 11457
rect 10170 11391 10566 11457
rect 16170 11391 16566 11457
rect 0 10978 800 11008
rect 18507 10978 19307 11008
rect 0 10918 2790 10978
rect 17496 10918 19307 10978
rect 0 10888 800 10918
rect 2730 10706 2790 10918
rect 4910 10847 5306 10913
rect 10910 10847 11306 10913
rect 16910 10847 17306 10913
rect 18507 10888 19307 10918
rect 2730 10646 11852 10706
rect 15840 10510 17050 10570
rect 0 10298 800 10328
rect 4170 10303 4566 10369
rect 10170 10303 10566 10369
rect 16170 10303 16566 10369
rect 16990 10298 17050 10510
rect 18507 10298 19307 10328
rect 0 10238 2790 10298
rect 16990 10238 19307 10298
rect 0 10208 800 10238
rect 2730 10162 2790 10238
rect 18507 10208 19307 10238
rect 2730 10102 9000 10162
rect 4910 9759 5306 9825
rect 10910 9759 11306 9825
rect 16910 9759 17306 9825
rect 0 9618 800 9648
rect 18507 9618 19307 9648
rect 0 9558 5504 9618
rect 17128 9558 19307 9618
rect 0 9528 800 9558
rect 18507 9528 19307 9558
rect 4170 9215 4566 9281
rect 10170 9215 10566 9281
rect 16170 9215 16566 9281
rect 0 8938 800 8968
rect 0 8878 1364 8938
rect 0 8848 800 8878
rect 4910 8671 5306 8737
rect 10910 8671 11306 8737
rect 16910 8671 17306 8737
rect 0 8258 800 8288
rect 0 8198 2790 8258
rect 0 8168 800 8198
rect 2730 7986 2790 8198
rect 4170 8127 4566 8193
rect 10170 8127 10566 8193
rect 16170 8127 16566 8193
rect 2730 7926 4768 7986
rect 2730 7790 7804 7850
rect 0 7578 800 7608
rect 2730 7578 2790 7790
rect 4910 7583 5306 7649
rect 10910 7583 11306 7649
rect 16910 7583 17306 7649
rect 0 7518 2790 7578
rect 0 7488 800 7518
rect 4170 7039 4566 7105
rect 10170 7039 10566 7105
rect 16170 7039 16566 7105
rect 0 6898 800 6928
rect 0 6838 10380 6898
rect 0 6808 800 6838
rect 4910 6495 5306 6561
rect 10910 6495 11306 6561
rect 16910 6495 17306 6561
rect 0 6218 800 6248
rect 0 6158 10380 6218
rect 0 6128 800 6158
rect 4170 5951 4566 6017
rect 10170 5951 10566 6017
rect 16170 5951 16566 6017
rect 0 5538 800 5568
rect 0 5478 2790 5538
rect 0 5448 800 5478
rect 2730 5266 2790 5478
rect 4910 5407 5306 5473
rect 10910 5407 11306 5473
rect 16910 5407 17306 5473
rect 2730 5206 8356 5266
rect 2730 5070 5964 5130
rect 0 4858 800 4888
rect 2730 4858 2790 5070
rect 4170 4863 4566 4929
rect 10170 4863 10566 4929
rect 16170 4863 16566 4929
rect 0 4798 2790 4858
rect 0 4768 800 4798
rect 4910 4319 5306 4385
rect 10910 4319 11306 4385
rect 16910 4319 17306 4385
rect 0 4178 800 4208
rect 0 4118 1364 4178
rect 0 4088 800 4118
rect 4170 3775 4566 3841
rect 10170 3775 10566 3841
rect 16170 3775 16566 3841
rect 0 3498 800 3528
rect 0 3438 4952 3498
rect 0 3408 800 3438
rect 4910 3231 5306 3297
rect 10910 3231 11306 3297
rect 16910 3231 17306 3297
rect 0 2818 800 2848
rect 0 2758 2192 2818
rect 0 2728 800 2758
rect 4170 2687 4566 2753
rect 10170 2687 10566 2753
rect 16170 2687 16566 2753
rect 4478 2350 6424 2410
rect 0 2138 800 2168
rect 4478 2138 4538 2350
rect 4910 2143 5306 2209
rect 10910 2143 11306 2209
rect 16910 2143 17306 2209
rect 0 2078 4538 2138
rect 0 2048 800 2078
rect 0 1458 800 1488
rect 0 1398 9000 1458
rect 0 1368 800 1398
rect 0 778 800 808
rect 0 718 12496 778
rect 0 688 800 718
rect 0 98 800 128
rect 0 38 12864 98
rect 0 8 800 38
<< metal4 >>
rect 4168 2128 4568 19088
rect 4908 2128 5308 19088
rect 10168 2128 10568 19088
rect 10908 2128 11308 19088
rect 16168 2128 16568 19088
rect 16908 2128 17308 19088
<< metal5 >>
rect 1056 18046 18172 18446
rect 1056 17306 18172 17706
rect 1056 12046 18172 12446
rect 1056 11306 18172 11706
rect 1056 6046 18172 6446
rect 1056 5306 18172 5706
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_0
timestamp 1571791925
transform 1 0 15364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_1
timestamp 1571791925
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_2
timestamp 1571791925
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_3
timestamp 1571791925
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_4
timestamp 1571791925
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_5
timestamp 1571791925
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_6
timestamp 1571791925
transform 1 0 16008 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_7
timestamp 1571791925
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_8
timestamp 1571791925
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_9
timestamp 1571791925
transform 1 0 14904 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_10
timestamp 1571791925
transform 1 0 16468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_11
timestamp 1571791925
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_12
timestamp 1571791925
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_13
timestamp 1571791925
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_14
timestamp 1571791925
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_15
timestamp 1571791925
transform 1 0 12052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_16
timestamp 1571791925
transform 1 0 14536 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_17
timestamp 1571791925
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_18
timestamp 1571791925
transform 1 0 15456 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_19
timestamp 1571791925
transform 1 0 14352 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_20
timestamp 1571791925
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_21
timestamp 1571791925
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_22
timestamp 1571791925
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_23
timestamp 1571791925
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_24
timestamp 1571791925
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_25
timestamp 1571791925
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_26
timestamp 1571791925
transform 1 0 13432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_27
timestamp 1571791925
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_28
timestamp 1571791925
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_29
timestamp 1571791925
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_30
timestamp 1571791925
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_31
timestamp 1571791925
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_32
timestamp 1571791925
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_33
timestamp 1571791925
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_34
timestamp 1571791925
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_35
timestamp 1571791925
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_36
timestamp 1571791925
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_37
timestamp 1571791925
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_38
timestamp 1571791925
transform 1 0 6808 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_39
timestamp 1571791925
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_40
timestamp 1571791925
transform 1 0 7636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_41
timestamp 1571791925
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_42
timestamp 1571791925
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_43
timestamp 1571791925
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_44
timestamp 1571791925
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_45
timestamp 1571791925
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_46
timestamp 1571791925
transform 1 0 6900 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_47
timestamp 1571791925
transform 1 0 4600 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_48
timestamp 1571791925
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_49
timestamp 1571791925
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_50
timestamp 1571791925
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_51
timestamp 1571791925
transform 1 0 16560 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_52
timestamp 1571791925
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_53
timestamp 1571791925
transform 1 0 15824 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_54
timestamp 1571791925
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_55
timestamp 1571791925
transform 1 0 11776 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_56
timestamp 1571791925
transform 1 0 11040 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_57
timestamp 1571791925
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_58
timestamp 1571791925
transform 1 0 12512 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_59
timestamp 1571791925
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_60
timestamp 1571791925
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_61
timestamp 1571791925
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_62
timestamp 1571791925
transform 1 0 15456 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_63
timestamp 1571791925
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_64
timestamp 1571791925
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_65
timestamp 1571791925
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_66
timestamp 1571791925
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_67
timestamp 1571791925
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_68
timestamp 1571791925
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_69
timestamp 1571791925
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_70
timestamp 1571791925
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_71
timestamp 1571791925
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_72
timestamp 1571791925
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_73
timestamp 1571791925
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_74
timestamp 1571791925
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_75
timestamp 1571791925
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_76
timestamp 1571791925
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_77
timestamp 1571791925
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_78
timestamp 1571791925
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_79
timestamp 1571791925
transform 1 0 14352 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_80
timestamp 1571791925
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_81
timestamp 1571791925
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_82
timestamp 1571791925
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_83
timestamp 1571791925
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_84
timestamp 1571791925
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_85
timestamp 1571791925
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_86
timestamp 1571791925
transform 1 0 9292 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_87
timestamp 1571791925
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_88
timestamp 1571791925
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_89
timestamp 1571791925
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_90
timestamp 1571791925
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_91
timestamp 1571791925
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_92
timestamp 1571791925
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_93
timestamp 1571791925
transform 1 0 9568 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_94
timestamp 1571791925
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  sky130_fd_sc_hd__a21o_2_0
timestamp 1571791925
transform -1 0 2300 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_0
timestamp 1571791925
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_1
timestamp 1571791925
transform 1 0 9936 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_2
timestamp 1571791925
transform 1 0 11040 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_3
timestamp 1571791925
transform -1 0 17296 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_4
timestamp 1571791925
transform 1 0 10212 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_5
timestamp 1571791925
transform 1 0 13248 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_6
timestamp 1571791925
transform 1 0 6532 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_7
timestamp 1571791925
transform 1 0 1932 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_8
timestamp 1571791925
transform 1 0 4232 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_9
timestamp 1571791925
transform 1 0 1472 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_10
timestamp 1571791925
transform 1 0 5704 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_11
timestamp 1571791925
transform 1 0 8004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_12
timestamp 1571791925
transform 1 0 5244 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_13
timestamp 1571791925
transform -1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_14
timestamp 1571791925
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_15
timestamp 1571791925
transform 1 0 5612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_16
timestamp 1571791925
transform 1 0 6992 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_17
timestamp 1571791925
transform 1 0 4508 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_18
timestamp 1571791925
transform 1 0 1748 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_19
timestamp 1571791925
transform 1 0 3404 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_20
timestamp 1571791925
transform 1 0 2484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_21
timestamp 1571791925
transform 1 0 5612 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_22
timestamp 1571791925
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_23
timestamp 1571791925
transform 1 0 16652 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_24
timestamp 1571791925
transform 1 0 12420 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_25
timestamp 1571791925
transform 1 0 10304 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_26
timestamp 1571791925
transform 1 0 11408 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_27
timestamp 1571791925
transform 1 0 14904 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_28
timestamp 1571791925
transform 1 0 9200 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_29
timestamp 1571791925
transform 1 0 1748 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  sky130_fd_sc_hd__a31o_2_30
timestamp 1571791925
transform 1 0 12972 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0
timestamp 1571791925
transform 1 0 15548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1571791925
transform -1 0 14904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_2
timestamp 1571791925
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_3
timestamp 1571791925
transform 1 0 10488 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_4
timestamp 1571791925
transform -1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_5
timestamp 1571791925
transform -1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_6
timestamp 1571791925
transform 1 0 12604 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_7
timestamp 1571791925
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_8
timestamp 1571791925
transform -1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_9
timestamp 1571791925
transform -1 0 3680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_10
timestamp 1571791925
transform 1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_11
timestamp 1571791925
transform -1 0 2944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_12
timestamp 1571791925
transform -1 0 9476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_13
timestamp 1571791925
transform -1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_14
timestamp 1571791925
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_15
timestamp 1571791925
transform -1 0 5888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_16
timestamp 1571791925
transform -1 0 5796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_17
timestamp 1571791925
transform -1 0 6808 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_18
timestamp 1571791925
transform -1 0 3588 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_19
timestamp 1571791925
transform -1 0 3220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_20
timestamp 1571791925
transform -1 0 4600 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_21
timestamp 1571791925
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_22
timestamp 1571791925
transform 1 0 8648 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_23
timestamp 1571791925
transform -1 0 6900 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_24
timestamp 1571791925
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_25
timestamp 1571791925
transform 1 0 17296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_26
timestamp 1571791925
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_27
timestamp 1571791925
transform -1 0 12696 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_28
timestamp 1571791925
transform -1 0 10212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_29
timestamp 1571791925
transform 1 0 11960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_30
timestamp 1571791925
transform -1 0 13984 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_31
timestamp 1571791925
transform 1 0 4508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0
timestamp 1571791925
transform -1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1571791925
transform 1 0 5152 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_2
timestamp 1571791925
transform 1 0 11408 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_3
timestamp 1571791925
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_0
timestamp 1571791925
transform 1 0 4876 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_1
timestamp 1571791925
transform 1 0 4600 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0
timestamp 1571791925
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1571791925
transform 1 0 11592 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_2
timestamp 1571791925
transform 1 0 5704 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_3
timestamp 1571791925
transform -1 0 6072 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_4
timestamp 1571791925
transform 1 0 4600 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_5
timestamp 1571791925
transform 1 0 5152 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_6
timestamp 1571791925
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_7
timestamp 1571791925
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_8
timestamp 1571791925
transform 1 0 8740 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1571791925
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1571791925
transform -1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1571791925
transform -1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1571791925
transform 1 0 14076 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1571791925
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1571791925
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1571791925
transform -1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1571791925
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1571791925
transform -1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1571791925
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1571791925
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1571791925
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1571791925
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1571791925
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1571791925
transform -1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1571791925
transform -1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1571791925
transform 1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1571791925
transform -1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1571791925
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1571791925
transform 1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1571791925
transform 1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1571791925
transform -1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1571791925
transform -1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1571791925
transform -1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1571791925
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1571791925
transform -1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1571791925
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1571791925
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1571791925
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1571791925
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1571791925
transform 1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1571791925
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1571791925
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1571791925
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1571791925
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1571791925
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1571791925
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_37
timestamp 1571791925
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_38
timestamp 1571791925
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_39
timestamp 1571791925
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_40
timestamp 1571791925
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_41
timestamp 1571791925
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_42
timestamp 1571791925
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_43
timestamp 1571791925
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_44
timestamp 1571791925
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_45
timestamp 1571791925
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_46
timestamp 1571791925
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_47
timestamp 1571791925
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_48
timestamp 1571791925
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_49
timestamp 1571791925
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_50
timestamp 1571791925
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_51
timestamp 1571791925
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_52
timestamp 1571791925
transform 1 0 7636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_53
timestamp 1571791925
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_54
timestamp 1571791925
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_55
timestamp 1571791925
transform 1 0 8004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_56
timestamp 1571791925
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_57
timestamp 1571791925
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_58
timestamp 1571791925
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_59
timestamp 1571791925
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_60
timestamp 1571791925
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_61
timestamp 1571791925
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_62
timestamp 1571791925
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_63
timestamp 1571791925
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_64
timestamp 1571791925
transform 1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_65
timestamp 1571791925
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_66
timestamp 1571791925
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_67
timestamp 1571791925
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_68
timestamp 1571791925
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_69
timestamp 1571791925
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_70
timestamp 1571791925
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_71
timestamp 1571791925
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_72
timestamp 1571791925
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_73
timestamp 1571791925
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_74
timestamp 1571791925
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_75
timestamp 1571791925
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_76
timestamp 1571791925
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_77
timestamp 1571791925
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_78
timestamp 1571791925
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_79
timestamp 1571791925
transform 1 0 4784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_80
timestamp 1571791925
transform 1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_81
timestamp 1571791925
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_82
timestamp 1571791925
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_83
timestamp 1571791925
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_84
timestamp 1571791925
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_85
timestamp 1571791925
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_86
timestamp 1571791925
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_87
timestamp 1571791925
transform -1 0 18124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_88
timestamp 1571791925
transform -1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_89
timestamp 1571791925
transform -1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_90
timestamp 1571791925
transform -1 0 18124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_91
timestamp 1571791925
transform -1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_92
timestamp 1571791925
transform -1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_93
timestamp 1571791925
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_94
timestamp 1571791925
transform 1 0 10212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_95
timestamp 1571791925
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_96
timestamp 1571791925
transform 1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_97
timestamp 1571791925
transform 1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_98
timestamp 1571791925
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_99
timestamp 1571791925
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_100
timestamp 1571791925
transform -1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_101
timestamp 1571791925
transform -1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_102
timestamp 1571791925
transform -1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_103
timestamp 1571791925
transform -1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_104
timestamp 1571791925
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_105
timestamp 1571791925
transform -1 0 18124 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_106
timestamp 1571791925
transform -1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_107
timestamp 1571791925
transform -1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_108
timestamp 1571791925
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_109
timestamp 1571791925
transform -1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_110
timestamp 1571791925
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_111
timestamp 1571791925
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_112
timestamp 1571791925
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_113
timestamp 1571791925
transform -1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_114
timestamp 1571791925
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1571791925
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1571791925
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1571791925
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1571791925
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1571791925
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1571791925
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1571791925
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1571791925
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1571791925
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1571791925
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_10
timestamp 1571791925
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_11
timestamp 1571791925
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_12
timestamp 1571791925
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_13
timestamp 1571791925
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_14
timestamp 1571791925
transform 1 0 4048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_15
timestamp 1571791925
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_16
timestamp 1571791925
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_17
timestamp 1571791925
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_18
timestamp 1571791925
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_19
timestamp 1571791925
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_20
timestamp 1571791925
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_21
timestamp 1571791925
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_22
timestamp 1571791925
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_23
timestamp 1571791925
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_24
timestamp 1571791925
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_25
timestamp 1571791925
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_26
timestamp 1571791925
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_27
timestamp 1571791925
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_28
timestamp 1571791925
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_29
timestamp 1571791925
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_30
timestamp 1571791925
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_31
timestamp 1571791925
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_32
timestamp 1571791925
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_33
timestamp 1571791925
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_34
timestamp 1571791925
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_35
timestamp 1571791925
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_36
timestamp 1571791925
transform 1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_37
timestamp 1571791925
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_38
timestamp 1571791925
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_39
timestamp 1571791925
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_40
timestamp 1571791925
transform 1 0 10396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_41
timestamp 1571791925
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_42
timestamp 1571791925
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_43
timestamp 1571791925
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_44
timestamp 1571791925
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_45
timestamp 1571791925
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_46
timestamp 1571791925
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_47
timestamp 1571791925
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_48
timestamp 1571791925
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_49
timestamp 1571791925
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_50
timestamp 1571791925
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1571791925
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1571791925
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1571791925
transform 1 0 17204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1571791925
transform 1 0 10120 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1571791925
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1571791925
transform 1 0 11684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1571791925
transform 1 0 17296 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1571791925
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1571791925
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1571791925
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1571791925
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1571791925
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1571791925
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1571791925
transform 1 0 3680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1571791925
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1571791925
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_16
timestamp 1571791925
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_17
timestamp 1571791925
transform 1 0 2392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_18
timestamp 1571791925
transform 1 0 4048 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_19
timestamp 1571791925
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_20
timestamp 1571791925
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_21
timestamp 1571791925
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_22
timestamp 1571791925
transform 1 0 6624 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_23
timestamp 1571791925
transform 1 0 7452 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_24
timestamp 1571791925
transform 1 0 5704 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_25
timestamp 1571791925
transform 1 0 6992 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_26
timestamp 1571791925
transform 1 0 6992 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_27
timestamp 1571791925
transform 1 0 4784 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_28
timestamp 1571791925
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_29
timestamp 1571791925
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_30
timestamp 1571791925
transform 1 0 9660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_31
timestamp 1571791925
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_32
timestamp 1571791925
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_33
timestamp 1571791925
transform 1 0 14720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1571791925
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1571791925
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1571791925
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1571791925
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1571791925
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1571791925
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1571791925
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1571791925
transform 1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1571791925
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1571791925
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1571791925
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1571791925
transform 1 0 13340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1571791925
transform 1 0 13432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1571791925
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1571791925
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1571791925
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1571791925
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1571791925
transform 1 0 2576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1571791925
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1571791925
transform 1 0 3404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1571791925
transform 1 0 6164 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1571791925
transform 1 0 7268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_22
timestamp 1571791925
transform 1 0 6900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_23
timestamp 1571791925
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_24
timestamp 1571791925
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_25
timestamp 1571791925
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_26
timestamp 1571791925
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_27
timestamp 1571791925
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_28
timestamp 1571791925
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_29
timestamp 1571791925
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_30
timestamp 1571791925
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_31
timestamp 1571791925
transform 1 0 4048 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_32
timestamp 1571791925
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_33
timestamp 1571791925
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_34
timestamp 1571791925
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_35
timestamp 1571791925
transform 1 0 16928 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_36
timestamp 1571791925
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_37
timestamp 1571791925
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_38
timestamp 1571791925
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_39
timestamp 1571791925
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_40
timestamp 1571791925
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_41
timestamp 1571791925
transform 1 0 10672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_42
timestamp 1571791925
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_43
timestamp 1571791925
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_44
timestamp 1571791925
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_45
timestamp 1571791925
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_46
timestamp 1571791925
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_47
timestamp 1571791925
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_48
timestamp 1571791925
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_49
timestamp 1571791925
transform 1 0 9476 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_0
timestamp 1571791925
transform 1 0 14076 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_1
timestamp 1571791925
transform 1 0 11316 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_2
timestamp 1571791925
transform -1 0 13708 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_3
timestamp 1571791925
transform 1 0 11040 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_4
timestamp 1571791925
transform 1 0 11500 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_5
timestamp 1571791925
transform 1 0 10672 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_6
timestamp 1571791925
transform -1 0 16008 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_7
timestamp 1571791925
transform 1 0 14444 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_8
timestamp 1571791925
transform 1 0 14628 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_9
timestamp 1571791925
transform 1 0 12788 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_10
timestamp 1571791925
transform 1 0 13616 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_11
timestamp 1571791925
transform -1 0 9476 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_12
timestamp 1571791925
transform 1 0 6164 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_13
timestamp 1571791925
transform -1 0 8280 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_14
timestamp 1571791925
transform 1 0 2024 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_15
timestamp 1571791925
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_16
timestamp 1571791925
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_17
timestamp 1571791925
transform 1 0 2852 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_18
timestamp 1571791925
transform 1 0 1748 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_19
timestamp 1571791925
transform 1 0 1380 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_20
timestamp 1571791925
transform -1 0 8648 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_21
timestamp 1571791925
transform 1 0 6348 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_22
timestamp 1571791925
transform -1 0 5704 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_23
timestamp 1571791925
transform 1 0 3956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_24
timestamp 1571791925
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_25
timestamp 1571791925
transform 1 0 4324 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_26
timestamp 1571791925
transform 1 0 4600 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_27
timestamp 1571791925
transform -1 0 8280 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_28
timestamp 1571791925
transform 1 0 6808 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_29
timestamp 1571791925
transform 1 0 2392 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_30
timestamp 1571791925
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_31
timestamp 1571791925
transform 1 0 1380 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_32
timestamp 1571791925
transform -1 0 3312 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_33
timestamp 1571791925
transform 1 0 3036 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_34
timestamp 1571791925
transform 1 0 1748 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_35
timestamp 1571791925
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_36
timestamp 1571791925
transform 1 0 6716 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_37
timestamp 1571791925
transform -1 0 9108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_38
timestamp 1571791925
transform -1 0 6624 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_39
timestamp 1571791925
transform 1 0 6624 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_40
timestamp 1571791925
transform 1 0 4324 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_41
timestamp 1571791925
transform 1 0 4324 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_42
timestamp 1571791925
transform 1 0 5060 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_43
timestamp 1571791925
transform 1 0 3772 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_44
timestamp 1571791925
transform 1 0 14628 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_45
timestamp 1571791925
transform 1 0 14076 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_46
timestamp 1571791925
transform 1 0 14444 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_47
timestamp 1571791925
transform -1 0 12420 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_48
timestamp 1571791925
transform 1 0 9660 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_49
timestamp 1571791925
transform 1 0 10212 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_50
timestamp 1571791925
transform 1 0 11500 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_51
timestamp 1571791925
transform 1 0 12880 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_52
timestamp 1571791925
transform 1 0 12972 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_53
timestamp 1571791925
transform 1 0 11960 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_54
timestamp 1571791925
transform -1 0 10856 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_55
timestamp 1571791925
transform 1 0 8280 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_56
timestamp 1571791925
transform 1 0 9384 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_57
timestamp 1571791925
transform 1 0 9476 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_58
timestamp 1571791925
transform 1 0 6348 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_59
timestamp 1571791925
transform 1 0 8004 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_60
timestamp 1571791925
transform 1 0 8188 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_61
timestamp 1571791925
transform -1 0 11040 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_62
timestamp 1571791925
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_63
timestamp 1571791925
transform 1 0 9108 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1571791925
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1571791925
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1571791925
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1571791925
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1571791925
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1571791925
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1571791925
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1571791925
transform 1 0 12696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1571791925
transform 1 0 11408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1571791925
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1571791925
transform 1 0 10120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1571791925
transform 1 0 12328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1571791925
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1571791925
transform 1 0 9752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1571791925
transform 1 0 9844 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1571791925
transform 1 0 10120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1571791925
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1571791925
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1571791925
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1571791925
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1571791925
transform 1 0 15364 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1571791925
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1571791925
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1571791925
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1571791925
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1571791925
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1571791925
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1571791925
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1571791925
transform 1 0 8096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1571791925
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1571791925
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1571791925
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1571791925
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1571791925
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1571791925
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1571791925
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1571791925
transform 1 0 4232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1571791925
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_38
timestamp 1571791925
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_39
timestamp 1571791925
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_40
timestamp 1571791925
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_41
timestamp 1571791925
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_42
timestamp 1571791925
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_43
timestamp 1571791925
transform 1 0 4416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_44
timestamp 1571791925
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_45
timestamp 1571791925
transform 1 0 4416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_46
timestamp 1571791925
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_47
timestamp 1571791925
transform 1 0 6900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_48
timestamp 1571791925
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_49
timestamp 1571791925
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_50
timestamp 1571791925
transform 1 0 8740 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_51
timestamp 1571791925
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_52
timestamp 1571791925
transform 1 0 5612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_53
timestamp 1571791925
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_54
timestamp 1571791925
transform 1 0 7636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_55
timestamp 1571791925
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_56
timestamp 1571791925
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_57
timestamp 1571791925
transform 1 0 2944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_58
timestamp 1571791925
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_59
timestamp 1571791925
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_60
timestamp 1571791925
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_61
timestamp 1571791925
transform 1 0 4968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_62
timestamp 1571791925
transform 1 0 2944 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_63
timestamp 1571791925
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_64
timestamp 1571791925
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_65
timestamp 1571791925
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_66
timestamp 1571791925
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_67
timestamp 1571791925
transform 1 0 8372 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_68
timestamp 1571791925
transform 1 0 7544 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_69
timestamp 1571791925
transform 1 0 7544 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_70
timestamp 1571791925
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_71
timestamp 1571791925
transform 1 0 15456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_72
timestamp 1571791925
transform 1 0 17756 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_73
timestamp 1571791925
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_74
timestamp 1571791925
transform 1 0 17756 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_75
timestamp 1571791925
transform 1 0 10120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_76
timestamp 1571791925
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_77
timestamp 1571791925
transform 1 0 10028 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_78
timestamp 1571791925
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_79
timestamp 1571791925
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_80
timestamp 1571791925
transform 1 0 10212 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_81
timestamp 1571791925
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_82
timestamp 1571791925
transform 1 0 17756 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_83
timestamp 1571791925
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_84
timestamp 1571791925
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_85
timestamp 1571791925
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_86
timestamp 1571791925
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_87
timestamp 1571791925
transform 1 0 17756 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_88
timestamp 1571791925
transform 1 0 11040 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_89
timestamp 1571791925
transform 1 0 14812 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_90
timestamp 1571791925
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_91
timestamp 1571791925
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_92
timestamp 1571791925
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_93
timestamp 1571791925
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_94
timestamp 1571791925
transform 1 0 15272 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_95
timestamp 1571791925
transform 1 0 10580 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_96
timestamp 1571791925
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_97
timestamp 1571791925
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_98
timestamp 1571791925
transform 1 0 9568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_99
timestamp 1571791925
transform 1 0 9568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0
timestamp 1571791925
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1571791925
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1571791925
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1571791925
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1571791925
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1571791925
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1571791925
transform 1 0 17664 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1571791925
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1571791925
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1571791925
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1571791925
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1571791925
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1571791925
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1571791925
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1571791925
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1571791925
transform 1 0 2208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1571791925
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1571791925
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1571791925
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1571791925
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1571791925
transform 1 0 6532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1571791925
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1571791925
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_23
timestamp 1571791925
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_24
timestamp 1571791925
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_25
timestamp 1571791925
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_26
timestamp 1571791925
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_27
timestamp 1571791925
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_28
timestamp 1571791925
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_29
timestamp 1571791925
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_30
timestamp 1571791925
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_31
timestamp 1571791925
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_32
timestamp 1571791925
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_33
timestamp 1571791925
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_34
timestamp 1571791925
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_35
timestamp 1571791925
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_36
timestamp 1571791925
transform 1 0 3128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_37
timestamp 1571791925
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_38
timestamp 1571791925
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_39
timestamp 1571791925
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_40
timestamp 1571791925
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_41
timestamp 1571791925
transform 1 0 12880 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_42
timestamp 1571791925
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_43
timestamp 1571791925
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_44
timestamp 1571791925
transform 1 0 17664 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_45
timestamp 1571791925
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_46
timestamp 1571791925
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_47
timestamp 1571791925
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1571791925
transform -1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1571791925
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1571791925
transform -1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1571791925
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1571791925
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1571791925
transform 1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1571791925
transform -1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1571791925
transform -1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1571791925
transform -1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1571791925
transform 1 0 12052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_10
timestamp 1571791925
transform -1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_11
timestamp 1571791925
transform 1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_12
timestamp 1571791925
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_13
timestamp 1571791925
transform 1 0 15364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_14
timestamp 1571791925
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_15
timestamp 1571791925
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_16
timestamp 1571791925
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_17
timestamp 1571791925
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_18
timestamp 1571791925
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_19
timestamp 1571791925
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_20
timestamp 1571791925
transform -1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_21
timestamp 1571791925
transform 1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_22
timestamp 1571791925
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_23
timestamp 1571791925
transform -1 0 5060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_24
timestamp 1571791925
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_25
timestamp 1571791925
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_26
timestamp 1571791925
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_27
timestamp 1571791925
transform -1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_28
timestamp 1571791925
transform -1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_29
timestamp 1571791925
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_30
timestamp 1571791925
transform 1 0 6992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_31
timestamp 1571791925
transform -1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_32
timestamp 1571791925
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_33
timestamp 1571791925
transform 1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_34
timestamp 1571791925
transform -1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_35
timestamp 1571791925
transform -1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_36
timestamp 1571791925
transform -1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_37
timestamp 1571791925
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_38
timestamp 1571791925
transform 1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_39
timestamp 1571791925
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_40
timestamp 1571791925
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_41
timestamp 1571791925
transform 1 0 1472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_42
timestamp 1571791925
transform -1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_43
timestamp 1571791925
transform -1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_44
timestamp 1571791925
transform -1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_45
timestamp 1571791925
transform 1 0 7636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_46
timestamp 1571791925
transform 1 0 7636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_47
timestamp 1571791925
transform -1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_48
timestamp 1571791925
transform -1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_49
timestamp 1571791925
transform -1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_50
timestamp 1571791925
transform -1 0 15180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_51
timestamp 1571791925
transform 1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_52
timestamp 1571791925
transform -1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_53
timestamp 1571791925
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_54
timestamp 1571791925
transform 1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_55
timestamp 1571791925
transform 1 0 12512 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_56
timestamp 1571791925
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_57
timestamp 1571791925
transform -1 0 10396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_58
timestamp 1571791925
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_59
timestamp 1571791925
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_60
timestamp 1571791925
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_61
timestamp 1571791925
transform -1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_62
timestamp 1571791925
transform 1 0 10672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_63
timestamp 1571791925
transform 1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_0
timestamp 1571791925
transform 1 0 12420 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_1
timestamp 1571791925
transform 1 0 10856 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_2
timestamp 1571791925
transform 1 0 12880 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_3
timestamp 1571791925
transform 1 0 10304 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_4
timestamp 1571791925
transform 1 0 17020 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_5
timestamp 1571791925
transform -1 0 17572 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_6
timestamp 1571791925
transform 1 0 6348 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_7
timestamp 1571791925
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_8
timestamp 1571791925
transform 1 0 7636 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_9
timestamp 1571791925
transform 1 0 1472 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_10
timestamp 1571791925
transform -1 0 4324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_11
timestamp 1571791925
transform 1 0 1748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_12
timestamp 1571791925
transform 1 0 8924 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_13
timestamp 1571791925
transform 1 0 7912 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_14
timestamp 1571791925
transform 1 0 5704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_15
timestamp 1571791925
transform 1 0 5888 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_16
timestamp 1571791925
transform 1 0 4876 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_17
timestamp 1571791925
transform 1 0 8832 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_18
timestamp 1571791925
transform 1 0 1380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_19
timestamp 1571791925
transform 1 0 4140 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_20
timestamp 1571791925
transform -1 0 2392 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_21
timestamp 1571791925
transform 1 0 4324 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_22
timestamp 1571791925
transform -1 0 7452 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_23
timestamp 1571791925
transform 1 0 2668 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_24
timestamp 1571791925
transform 1 0 5336 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_25
timestamp 1571791925
transform -1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_26
timestamp 1571791925
transform 1 0 10948 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_27
timestamp 1571791925
transform 1 0 11776 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_28
timestamp 1571791925
transform 1 0 12696 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_29
timestamp 1571791925
transform 1 0 10948 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_30
timestamp 1571791925
transform 1 0 9200 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  sky130_fd_sc_hd__nand3_2_0
timestamp 1571791925
transform -1 0 2576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1571791925
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1571791925
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1571791925
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1571791925
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1571791925
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1571791925
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1571791925
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1571791925
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1571791925
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1571791925
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1571791925
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1571791925
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1571791925
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1571791925
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1571791925
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1571791925
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1571791925
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1571791925
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1571791925
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1571791925
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1571791925
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1571791925
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1571791925
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1571791925
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1571791925
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1571791925
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1571791925
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1571791925
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1571791925
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1571791925
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1571791925
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1571791925
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1571791925
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1571791925
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1571791925
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1571791925
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1571791925
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1571791925
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1571791925
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1571791925
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1571791925
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1571791925
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1571791925
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1571791925
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1571791925
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1571791925
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1571791925
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1571791925
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1571791925
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1571791925
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1571791925
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1571791925
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1571791925
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1571791925
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1571791925
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1571791925
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1571791925
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1571791925
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1571791925
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1571791925
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1571791925
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1571791925
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1571791925
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1571791925
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1571791925
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1571791925
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1571791925
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1571791925
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1571791925
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1571791925
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1571791925
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1571791925
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1571791925
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1571791925
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1571791925
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1571791925
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1571791925
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1571791925
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1571791925
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1571791925
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1571791925
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1571791925
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1571791925
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1571791925
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1571791925
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1571791925
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1571791925
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1571791925
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1571791925
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1571791925
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1571791925
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1571791925
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1571791925
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1571791925
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1571791925
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1571791925
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1571791925
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1571791925
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1571791925
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_0
timestamp 1571791925
transform -1 0 13432 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_1
timestamp 1571791925
transform -1 0 12696 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_2
timestamp 1571791925
transform 1 0 10212 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_3
timestamp 1571791925
transform -1 0 17848 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_4
timestamp 1571791925
transform 1 0 12788 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_5
timestamp 1571791925
transform 1 0 7544 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_6
timestamp 1571791925
transform 1 0 6348 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_7
timestamp 1571791925
transform -1 0 5244 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_8
timestamp 1571791925
transform 1 0 1656 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_9
timestamp 1571791925
transform 1 0 3680 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_10
timestamp 1571791925
transform -1 0 7544 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_11
timestamp 1571791925
transform -1 0 9016 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_12
timestamp 1571791925
transform 1 0 1564 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_13
timestamp 1571791925
transform 1 0 6440 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_14
timestamp 1571791925
transform 1 0 1840 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_15
timestamp 1571791925
transform 1 0 1748 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_16
timestamp 1571791925
transform 1 0 3956 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_17
timestamp 1571791925
transform 1 0 5796 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_18
timestamp 1571791925
transform 1 0 4416 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_19
timestamp 1571791925
transform -1 0 2668 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_20
timestamp 1571791925
transform -1 0 15824 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_21
timestamp 1571791925
transform -1 0 12696 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_22
timestamp 1571791925
transform 1 0 12236 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_23
timestamp 1571791925
transform 1 0 10764 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_24
timestamp 1571791925
transform 1 0 12052 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_25
timestamp 1571791925
transform -1 0 10120 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_26
timestamp 1571791925
transform 1 0 8464 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_27
timestamp 1571791925
transform 1 0 5060 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_28
timestamp 1571791925
transform -1 0 17848 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_29
timestamp 1571791925
transform 1 0 8924 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  sky130_fd_sc_hd__xnor2_2_30
timestamp 1571791925
transform 1 0 8924 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_0
timestamp 1571791925
transform -1 0 15364 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_1
timestamp 1571791925
transform -1 0 15824 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_2
timestamp 1571791925
transform -1 0 11776 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_3
timestamp 1571791925
transform 1 0 10212 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_4
timestamp 1571791925
transform -1 0 13432 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_5
timestamp 1571791925
transform -1 0 11132 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_6
timestamp 1571791925
transform 1 0 16376 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_7
timestamp 1571791925
transform 1 0 6348 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_8
timestamp 1571791925
transform -1 0 8556 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_9
timestamp 1571791925
transform -1 0 4968 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_10
timestamp 1571791925
transform -1 0 3312 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_11
timestamp 1571791925
transform 1 0 6348 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_12
timestamp 1571791925
transform -1 0 8832 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_13
timestamp 1571791925
transform -1 0 5336 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_14
timestamp 1571791925
transform 1 0 4508 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_15
timestamp 1571791925
transform -1 0 8832 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_16
timestamp 1571791925
transform 1 0 8096 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_17
timestamp 1571791925
transform 1 0 6440 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_18
timestamp 1571791925
transform -1 0 4048 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_19
timestamp 1571791925
transform -1 0 4968 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_20
timestamp 1571791925
transform 1 0 3128 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_21
timestamp 1571791925
transform 1 0 7636 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_22
timestamp 1571791925
transform -1 0 6256 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_23
timestamp 1571791925
transform -1 0 16008 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_24
timestamp 1571791925
transform 1 0 16376 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_25
timestamp 1571791925
transform -1 0 11408 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_26
timestamp 1571791925
transform -1 0 14536 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_27
timestamp 1571791925
transform -1 0 12880 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_28
timestamp 1571791925
transform -1 0 10764 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_29
timestamp 1571791925
transform 1 0 11776 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  sky130_fd_sc_hd__xor2_2_30
timestamp 1571791925
transform -1 0 3588 0 -1 10880
box -38 -48 1234 592
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_0
timestamp 1571791925
transform 1 0 15410 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_1
timestamp 1571791925
transform 1 0 14306 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_2
timestamp 1571791925
transform 1 0 15594 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_3
timestamp 1571791925
transform 1 0 14858 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_4
timestamp 1571791925
transform 1 0 14858 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_5
timestamp 1571791925
transform 1 0 13938 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_6
timestamp 1571791925
transform 1 0 14214 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_7
timestamp 1571791925
transform 1 0 15502 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_8
timestamp 1571791925
transform 1 0 14398 0 1 4522
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_9
timestamp 1571791925
transform 1 0 13662 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_10
timestamp 1571791925
transform 1 0 14950 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_11
timestamp 1571791925
transform 1 0 13938 0 1 4522
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_12
timestamp 1571791925
transform 1 0 14122 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_13
timestamp 1571791925
transform 1 0 13662 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_14
timestamp 1571791925
transform 1 0 14674 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_15
timestamp 1571791925
transform 1 0 14490 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_16
timestamp 1571791925
transform 1 0 15962 0 1 3162
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_17
timestamp 1571791925
transform 1 0 15778 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_18
timestamp 1571791925
transform 1 0 15870 0 1 4454
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_19
timestamp 1571791925
transform 1 0 14674 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_20
timestamp 1571791925
transform 1 0 14950 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_21
timestamp 1571791925
transform 1 0 14858 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_22
timestamp 1571791925
transform 1 0 14398 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_23
timestamp 1571791925
transform 1 0 14674 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_24
timestamp 1571791925
transform 1 0 13018 0 1 2618
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_25
timestamp 1571791925
transform 1 0 12466 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_26
timestamp 1571791925
transform 1 0 12834 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_27
timestamp 1571791925
transform 1 0 12742 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_28
timestamp 1571791925
transform 1 0 13110 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_29
timestamp 1571791925
transform 1 0 9706 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_30
timestamp 1571791925
transform 1 0 9982 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_31
timestamp 1571791925
transform 1 0 10718 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_32
timestamp 1571791925
transform 1 0 10166 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_33
timestamp 1571791925
transform 1 0 10258 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_34
timestamp 1571791925
transform 1 0 10626 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_35
timestamp 1571791925
transform 1 0 10994 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_36
timestamp 1571791925
transform 1 0 9982 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_37
timestamp 1571791925
transform 1 0 10902 0 1 3910
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_38
timestamp 1571791925
transform 1 0 10902 0 1 4794
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_39
timestamp 1571791925
transform 1 0 10534 0 1 4658
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_40
timestamp 1571791925
transform 1 0 9614 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_41
timestamp 1571791925
transform 1 0 9982 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_42
timestamp 1571791925
transform 1 0 9798 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_43
timestamp 1571791925
transform 1 0 10074 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_44
timestamp 1571791925
transform 1 0 10534 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_45
timestamp 1571791925
transform 1 0 10350 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_46
timestamp 1571791925
transform 1 0 10534 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_47
timestamp 1571791925
transform 1 0 9890 0 1 4794
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_48
timestamp 1571791925
transform 1 0 11270 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_49
timestamp 1571791925
transform 1 0 11362 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_50
timestamp 1571791925
transform 1 0 11914 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_51
timestamp 1571791925
transform 1 0 13294 0 1 4182
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_52
timestamp 1571791925
transform 1 0 12926 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_53
timestamp 1571791925
transform 1 0 13294 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_54
timestamp 1571791925
transform 1 0 13478 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_55
timestamp 1571791925
transform 1 0 13018 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_56
timestamp 1571791925
transform 1 0 11914 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_57
timestamp 1571791925
transform 1 0 11638 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_58
timestamp 1571791925
transform 1 0 13386 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_59
timestamp 1571791925
transform 1 0 12282 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_60
timestamp 1571791925
transform 1 0 11638 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_61
timestamp 1571791925
transform 1 0 13202 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_62
timestamp 1571791925
transform 1 0 13294 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_63
timestamp 1571791925
transform 1 0 11638 0 1 4658
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_64
timestamp 1571791925
transform 1 0 11730 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_65
timestamp 1571791925
transform 1 0 12282 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_66
timestamp 1571791925
transform 1 0 11914 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_67
timestamp 1571791925
transform 1 0 11546 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_68
timestamp 1571791925
transform 1 0 13110 0 1 6222
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_69
timestamp 1571791925
transform 1 0 12282 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_70
timestamp 1571791925
transform 1 0 11638 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_71
timestamp 1571791925
transform 1 0 12742 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_72
timestamp 1571791925
transform 1 0 12558 0 1 7718
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_73
timestamp 1571791925
transform 1 0 12374 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_74
timestamp 1571791925
transform 1 0 12834 0 1 6222
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_75
timestamp 1571791925
transform 1 0 13110 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_76
timestamp 1571791925
transform 1 0 12098 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_77
timestamp 1571791925
transform 1 0 12190 0 1 7718
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_78
timestamp 1571791925
transform 1 0 13478 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_79
timestamp 1571791925
transform 1 0 11638 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_80
timestamp 1571791925
transform 1 0 13570 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_81
timestamp 1571791925
transform 1 0 12466 0 1 6086
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_82
timestamp 1571791925
transform 1 0 13294 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_83
timestamp 1571791925
transform 1 0 11914 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_84
timestamp 1571791925
transform 1 0 11822 0 1 7310
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_85
timestamp 1571791925
transform 1 0 12926 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_86
timestamp 1571791925
transform 1 0 13294 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_87
timestamp 1571791925
transform 1 0 13294 0 1 5814
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_88
timestamp 1571791925
transform 1 0 10810 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_89
timestamp 1571791925
transform 1 0 10074 0 1 7446
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_90
timestamp 1571791925
transform 1 0 11362 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_91
timestamp 1571791925
transform 1 0 11270 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_92
timestamp 1571791925
transform 1 0 11362 0 1 5746
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_93
timestamp 1571791925
transform 1 0 9798 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_94
timestamp 1571791925
transform 1 0 10994 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_95
timestamp 1571791925
transform 1 0 10626 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_96
timestamp 1571791925
transform 1 0 10810 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_97
timestamp 1571791925
transform 1 0 10626 0 1 6426
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_98
timestamp 1571791925
transform 1 0 10442 0 1 6358
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_99
timestamp 1571791925
transform 1 0 11178 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_100
timestamp 1571791925
transform 1 0 11454 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_101
timestamp 1571791925
transform 1 0 10718 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_102
timestamp 1571791925
transform 1 0 10902 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_103
timestamp 1571791925
transform 1 0 10554 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_104
timestamp 1571791925
transform 1 0 11362 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_105
timestamp 1571791925
transform 1 0 10166 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_106
timestamp 1571791925
transform 1 0 10350 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_107
timestamp 1571791925
transform 1 0 11270 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_108
timestamp 1571791925
transform 1 0 11086 0 1 6902
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_109
timestamp 1571791925
transform 1 0 10534 0 1 5746
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_110
timestamp 1571791925
transform 1 0 10718 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_111
timestamp 1571791925
transform 1 0 10258 0 1 6154
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_112
timestamp 1571791925
transform 1 0 10994 0 1 10098
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_113
timestamp 1571791925
transform 1 0 11362 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_114
timestamp 1571791925
transform 1 0 10534 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_115
timestamp 1571791925
transform 1 0 9614 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_116
timestamp 1571791925
transform 1 0 10534 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_117
timestamp 1571791925
transform 1 0 9982 0 1 10098
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_118
timestamp 1571791925
transform 1 0 9798 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_119
timestamp 1571791925
transform 1 0 11086 0 1 9010
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_120
timestamp 1571791925
transform 1 0 10718 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_121
timestamp 1571791925
transform 1 0 10350 0 1 9350
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_122
timestamp 1571791925
transform 1 0 9982 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_123
timestamp 1571791925
transform 1 0 9982 0 1 9350
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_124
timestamp 1571791925
transform 1 0 10810 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_125
timestamp 1571791925
transform 1 0 9890 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_126
timestamp 1571791925
transform 1 0 10718 0 1 9486
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_127
timestamp 1571791925
transform 1 0 10718 0 1 9146
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_128
timestamp 1571791925
transform 1 0 13018 0 1 10506
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_129
timestamp 1571791925
transform 1 0 12650 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_130
timestamp 1571791925
transform 1 0 12466 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_131
timestamp 1571791925
transform 1 0 12006 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_132
timestamp 1571791925
transform 1 0 13018 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_133
timestamp 1571791925
transform 1 0 12098 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_134
timestamp 1571791925
transform 1 0 12834 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_135
timestamp 1571791925
transform 1 0 13202 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_136
timestamp 1571791925
transform 1 0 12834 0 1 8806
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_137
timestamp 1571791925
transform 1 0 11638 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_138
timestamp 1571791925
transform 1 0 13110 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_139
timestamp 1571791925
transform 1 0 13386 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_140
timestamp 1571791925
transform 1 0 11914 0 1 9622
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_141
timestamp 1571791925
transform 1 0 11546 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_142
timestamp 1571791925
transform 1 0 17066 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_143
timestamp 1571791925
transform 1 0 17342 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_144
timestamp 1571791925
transform 1 0 17434 0 1 7922
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_145
timestamp 1571791925
transform 1 0 15962 0 1 7922
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_146
timestamp 1571791925
transform 1 0 13662 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_147
timestamp 1571791925
transform 1 0 14398 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_148
timestamp 1571791925
transform 1 0 14214 0 1 7718
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_149
timestamp 1571791925
transform 1 0 14214 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_150
timestamp 1571791925
transform 1 0 14306 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_151
timestamp 1571791925
transform 1 0 14306 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_152
timestamp 1571791925
transform 1 0 14214 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_153
timestamp 1571791925
transform 1 0 13846 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_154
timestamp 1571791925
transform 1 0 14582 0 1 6086
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_155
timestamp 1571791925
transform 1 0 15042 0 1 5746
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_156
timestamp 1571791925
transform 1 0 15410 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_157
timestamp 1571791925
transform 1 0 15502 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_158
timestamp 1571791925
transform 1 0 14766 0 1 9010
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_159
timestamp 1571791925
transform 1 0 14490 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_160
timestamp 1571791925
transform 1 0 14674 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_161
timestamp 1571791925
transform 1 0 15594 0 1 9622
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_162
timestamp 1571791925
transform 1 0 15502 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_163
timestamp 1571791925
transform 1 0 14950 0 1 10098
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_164
timestamp 1571791925
transform 1 0 16422 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_165
timestamp 1571791925
transform 1 0 16698 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_166
timestamp 1571791925
transform 1 0 17434 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_167
timestamp 1571791925
transform 1 0 17526 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_168
timestamp 1571791925
transform 1 0 17526 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_169
timestamp 1571791925
transform 1 0 17066 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_170
timestamp 1571791925
transform 1 0 17342 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_171
timestamp 1571791925
transform 1 0 17434 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_172
timestamp 1571791925
transform 1 0 17250 0 1 9418
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_173
timestamp 1571791925
transform 1 0 17526 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_174
timestamp 1571791925
transform 1 0 16974 0 1 9690
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_175
timestamp 1571791925
transform 1 0 16698 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_176
timestamp 1571791925
transform 1 0 16238 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_177
timestamp 1571791925
transform 1 0 16422 0 1 9894
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_178
timestamp 1571791925
transform 1 0 16146 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_179
timestamp 1571791925
transform 1 0 16514 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_180
timestamp 1571791925
transform 1 0 16238 0 1 9010
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_181
timestamp 1571791925
transform 1 0 16698 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_182
timestamp 1571791925
transform 1 0 17342 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_183
timestamp 1571791925
transform 1 0 16882 0 1 9690
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_184
timestamp 1571791925
transform 1 0 15686 0 1 7786
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_185
timestamp 1571791925
transform 1 0 12834 0 1 5338
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_186
timestamp 1571791925
transform 1 0 14490 0 1 5338
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_187
timestamp 1571791925
transform 1 0 7682 0 1 2618
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_188
timestamp 1571791925
transform 1 0 7866 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_189
timestamp 1571791925
transform 1 0 8050 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_190
timestamp 1571791925
transform 1 0 9062 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_191
timestamp 1571791925
transform 1 0 6394 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_192
timestamp 1571791925
transform 1 0 7222 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_193
timestamp 1571791925
transform 1 0 6670 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_194
timestamp 1571791925
transform 1 0 6762 0 1 2482
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_195
timestamp 1571791925
transform 1 0 7314 0 1 2618
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_196
timestamp 1571791925
transform 1 0 6486 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_197
timestamp 1571791925
transform 1 0 5750 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_198
timestamp 1571791925
transform 1 0 6578 0 1 3978
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_199
timestamp 1571791925
transform 1 0 6118 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_200
timestamp 1571791925
transform 1 0 6210 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_201
timestamp 1571791925
transform 1 0 7130 0 1 4182
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_202
timestamp 1571791925
transform 1 0 5750 0 1 4658
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_203
timestamp 1571791925
transform 1 0 5842 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_204
timestamp 1571791925
transform 1 0 6302 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_205
timestamp 1571791925
transform 1 0 7406 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_206
timestamp 1571791925
transform 1 0 6946 0 1 4250
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_207
timestamp 1571791925
transform 1 0 5566 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_208
timestamp 1571791925
transform 1 0 5658 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_209
timestamp 1571791925
transform 1 0 7406 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_210
timestamp 1571791925
transform 1 0 5474 0 1 3706
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_211
timestamp 1571791925
transform 1 0 6210 0 1 4794
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_212
timestamp 1571791925
transform 1 0 6486 0 1 4726
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_213
timestamp 1571791925
transform 1 0 6854 0 1 4250
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_214
timestamp 1571791925
transform 1 0 6762 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_215
timestamp 1571791925
transform 1 0 6762 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_216
timestamp 1571791925
transform 1 0 6946 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_217
timestamp 1571791925
transform 1 0 6026 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_218
timestamp 1571791925
transform 1 0 6118 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_219
timestamp 1571791925
transform 1 0 6670 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_220
timestamp 1571791925
transform 1 0 9430 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_221
timestamp 1571791925
transform 1 0 7682 0 1 3162
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_222
timestamp 1571791925
transform 1 0 9062 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_223
timestamp 1571791925
transform 1 0 8234 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_224
timestamp 1571791925
transform 1 0 7958 0 1 3706
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_225
timestamp 1571791925
transform 1 0 8234 0 1 4046
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_226
timestamp 1571791925
transform 1 0 7682 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_227
timestamp 1571791925
transform 1 0 9154 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_228
timestamp 1571791925
transform 1 0 9246 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_229
timestamp 1571791925
transform 1 0 8510 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_230
timestamp 1571791925
transform 1 0 7866 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_231
timestamp 1571791925
transform 1 0 9246 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_232
timestamp 1571791925
transform 1 0 9338 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_233
timestamp 1571791925
transform 1 0 8050 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_234
timestamp 1571791925
transform 1 0 9338 0 1 4794
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_235
timestamp 1571791925
transform 1 0 7958 0 1 4522
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_236
timestamp 1571791925
transform 1 0 7498 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_237
timestamp 1571791925
transform 1 0 8234 0 1 4658
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_238
timestamp 1571791925
transform 1 0 3542 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_239
timestamp 1571791925
transform 1 0 3450 0 1 2618
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_240
timestamp 1571791925
transform 1 0 2530 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_241
timestamp 1571791925
transform 1 0 1978 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_242
timestamp 1571791925
transform 1 0 2438 0 1 2618
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_243
timestamp 1571791925
transform 1 0 2162 0 1 2414
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_244
timestamp 1571791925
transform 1 0 3266 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_245
timestamp 1571791925
transform 1 0 1794 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_246
timestamp 1571791925
transform 1 0 1702 0 1 4182
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_247
timestamp 1571791925
transform 1 0 2162 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_248
timestamp 1571791925
transform 1 0 2530 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_249
timestamp 1571791925
transform 1 0 1702 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_250
timestamp 1571791925
transform 1 0 3174 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_251
timestamp 1571791925
transform 1 0 2070 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_252
timestamp 1571791925
transform 1 0 2346 0 1 4046
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_253
timestamp 1571791925
transform 1 0 1426 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_254
timestamp 1571791925
transform 1 0 2530 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_255
timestamp 1571791925
transform 1 0 1886 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_256
timestamp 1571791925
transform 1 0 2622 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_257
timestamp 1571791925
transform 1 0 2346 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_258
timestamp 1571791925
transform 1 0 2714 0 1 3910
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_259
timestamp 1571791925
transform 1 0 2162 0 1 3910
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_260
timestamp 1571791925
transform 1 0 1518 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_261
timestamp 1571791925
transform 1 0 1794 0 1 4182
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_262
timestamp 1571791925
transform 1 0 1978 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_263
timestamp 1571791925
transform 1 0 1978 0 1 5270
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_264
timestamp 1571791925
transform 1 0 4278 0 1 3978
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_265
timestamp 1571791925
transform 1 0 4002 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_266
timestamp 1571791925
transform 1 0 3542 0 1 3502
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_267
timestamp 1571791925
transform 1 0 4830 0 1 4182
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_268
timestamp 1571791925
transform 1 0 4830 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_269
timestamp 1571791925
transform 1 0 3450 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_270
timestamp 1571791925
transform 1 0 5014 0 1 3978
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_271
timestamp 1571791925
transform 1 0 4278 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_272
timestamp 1571791925
transform 1 0 4646 0 1 4590
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_273
timestamp 1571791925
transform 1 0 4462 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_274
timestamp 1571791925
transform 1 0 3634 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_275
timestamp 1571791925
transform 1 0 5198 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_276
timestamp 1571791925
transform 1 0 4600 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_277
timestamp 1571791925
transform 1 0 4922 0 1 4114
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_278
timestamp 1571791925
transform 1 0 3450 0 1 3434
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_279
timestamp 1571791925
transform 1 0 4278 0 1 3094
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_280
timestamp 1571791925
transform 1 0 4370 0 1 5202
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_281
timestamp 1571791925
transform 1 0 3818 0 1 2958
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_282
timestamp 1571791925
transform 1 0 5014 0 1 3570
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_283
timestamp 1571791925
transform 1 0 4646 0 1 5134
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_284
timestamp 1571791925
transform 1 0 4646 0 1 4250
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_285
timestamp 1571791925
transform 1 0 4186 0 1 4658
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_286
timestamp 1571791925
transform 1 0 5290 0 1 6698
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_287
timestamp 1571791925
transform 1 0 4922 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_288
timestamp 1571791925
transform 1 0 5014 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_289
timestamp 1571791925
transform 1 0 3542 0 1 6970
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_290
timestamp 1571791925
transform 1 0 5290 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_291
timestamp 1571791925
transform 1 0 4002 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_292
timestamp 1571791925
transform 1 0 4278 0 1 6358
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_293
timestamp 1571791925
transform 1 0 4554 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_294
timestamp 1571791925
transform 1 0 4554 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_295
timestamp 1571791925
transform 1 0 4002 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_296
timestamp 1571791925
transform 1 0 3910 0 1 6698
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_297
timestamp 1571791925
transform 1 0 3818 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_298
timestamp 1571791925
transform 1 0 4646 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_299
timestamp 1571791925
transform 1 0 4830 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_300
timestamp 1571791925
transform 1 0 1886 0 1 5610
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_301
timestamp 1571791925
transform 1 0 2162 0 1 6222
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_302
timestamp 1571791925
transform 1 0 2162 0 1 7514
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_303
timestamp 1571791925
transform 1 0 1702 0 1 7922
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_304
timestamp 1571791925
transform 1 0 1426 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_305
timestamp 1571791925
transform 1 0 2070 0 1 6698
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_306
timestamp 1571791925
transform 1 0 1610 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_307
timestamp 1571791925
transform 1 0 2714 0 1 6426
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_308
timestamp 1571791925
transform 1 0 1794 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_309
timestamp 1571791925
transform 1 0 2070 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_310
timestamp 1571791925
transform 1 0 1886 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_311
timestamp 1571791925
transform 1 0 1794 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_312
timestamp 1571791925
transform 1 0 1794 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_313
timestamp 1571791925
transform 1 0 2162 0 1 9486
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_314
timestamp 1571791925
transform 1 0 3174 0 1 9622
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_315
timestamp 1571791925
transform 1 0 2898 0 1 9486
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_316
timestamp 1571791925
transform 1 0 2898 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_317
timestamp 1571791925
transform 1 0 2806 0 1 9622
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_318
timestamp 1571791925
transform 1 0 2070 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_319
timestamp 1571791925
transform 1 0 2530 0 1 8806
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_320
timestamp 1571791925
transform 1 0 1886 0 1 9146
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_321
timestamp 1571791925
transform 1 0 1886 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_322
timestamp 1571791925
transform 1 0 1978 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_323
timestamp 1571791925
transform 1 0 2070 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_324
timestamp 1571791925
transform 1 0 1518 0 1 8330
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_325
timestamp 1571791925
transform 1 0 2714 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_326
timestamp 1571791925
transform 1 0 2990 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_327
timestamp 1571791925
transform 1 0 3266 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_328
timestamp 1571791925
transform 1 0 2162 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_329
timestamp 1571791925
transform 1 0 1702 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_330
timestamp 1571791925
transform 1 0 3174 0 1 8058
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_331
timestamp 1571791925
transform 1 0 4830 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_332
timestamp 1571791925
transform 1 0 3910 0 1 9894
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_333
timestamp 1571791925
transform 1 0 4922 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_334
timestamp 1571791925
transform 1 0 3910 0 1 8058
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_335
timestamp 1571791925
transform 1 0 4646 0 1 9010
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_336
timestamp 1571791925
transform 1 0 4922 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_337
timestamp 1571791925
transform 1 0 4002 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_338
timestamp 1571791925
transform 1 0 3910 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_339
timestamp 1571791925
transform 1 0 4462 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_340
timestamp 1571791925
transform 1 0 3818 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_341
timestamp 1571791925
transform 1 0 4646 0 1 9690
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_342
timestamp 1571791925
transform 1 0 4278 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_343
timestamp 1571791925
transform 1 0 4830 0 1 10098
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_344
timestamp 1571791925
transform 1 0 4094 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_345
timestamp 1571791925
transform 1 0 4554 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_346
timestamp 1571791925
transform 1 0 3358 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_347
timestamp 1571791925
transform 1 0 8694 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_348
timestamp 1571791925
transform 1 0 8142 0 1 6426
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_349
timestamp 1571791925
transform 1 0 9062 0 1 5542
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_350
timestamp 1571791925
transform 1 0 7590 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_351
timestamp 1571791925
transform 1 0 8326 0 1 7310
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_352
timestamp 1571791925
transform 1 0 7774 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_353
timestamp 1571791925
transform 1 0 7958 0 1 5746
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_354
timestamp 1571791925
transform 1 0 7498 0 1 6086
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_355
timestamp 1571791925
transform 1 0 8346 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_356
timestamp 1571791925
transform 1 0 9246 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_357
timestamp 1571791925
transform 1 0 8602 0 1 6358
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_358
timestamp 1571791925
transform 1 0 8142 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_359
timestamp 1571791925
transform 1 0 9062 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_360
timestamp 1571791925
transform 1 0 8050 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_361
timestamp 1571791925
transform 1 0 8050 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_362
timestamp 1571791925
transform 1 0 7682 0 1 7174
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_363
timestamp 1571791925
transform 1 0 9338 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_364
timestamp 1571791925
transform 1 0 8234 0 1 6290
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_365
timestamp 1571791925
transform 1 0 8418 0 1 6426
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_366
timestamp 1571791925
transform 1 0 8694 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_367
timestamp 1571791925
transform 1 0 7958 0 1 7786
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_368
timestamp 1571791925
transform 1 0 5658 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_369
timestamp 1571791925
transform 1 0 6118 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_370
timestamp 1571791925
transform 1 0 5566 0 1 6630
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_371
timestamp 1571791925
transform 1 0 5842 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_372
timestamp 1571791925
transform 1 0 6302 0 1 6834
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_373
timestamp 1571791925
transform 1 0 5934 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_374
timestamp 1571791925
transform 1 0 6026 0 1 7718
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_375
timestamp 1571791925
transform 1 0 5658 0 1 7922
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_376
timestamp 1571791925
transform 1 0 7038 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_377
timestamp 1571791925
transform 1 0 5750 0 1 5678
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_378
timestamp 1571791925
transform 1 0 6394 0 1 6766
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_379
timestamp 1571791925
transform 1 0 7038 0 1 5814
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_380
timestamp 1571791925
transform 1 0 6026 0 1 7446
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_381
timestamp 1571791925
transform 1 0 6302 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_382
timestamp 1571791925
transform 1 0 7406 0 1 7378
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_383
timestamp 1571791925
transform 1 0 5934 0 1 7854
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_384
timestamp 1571791925
transform 1 0 5474 0 1 6698
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_385
timestamp 1571791925
transform 1 0 6118 0 1 7718
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_386
timestamp 1571791925
transform 1 0 5750 0 1 6086
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_387
timestamp 1571791925
transform 1 0 6486 0 1 7310
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_388
timestamp 1571791925
transform 1 0 6651 0 1 6970
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_389
timestamp 1571791925
transform 1 0 5750 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_390
timestamp 1571791925
transform 1 0 7130 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_391
timestamp 1571791925
transform 1 0 6486 0 1 9350
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_392
timestamp 1571791925
transform 1 0 7222 0 1 8534
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_393
timestamp 1571791925
transform 1 0 6394 0 1 9146
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_394
timestamp 1571791925
transform 1 0 5750 0 1 7990
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_395
timestamp 1571791925
transform 1 0 6026 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_396
timestamp 1571791925
transform 1 0 6486 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_397
timestamp 1571791925
transform 1 0 6670 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_398
timestamp 1571791925
transform 1 0 6118 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_399
timestamp 1571791925
transform 1 0 6210 0 1 10574
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_400
timestamp 1571791925
transform 1 0 7038 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_401
timestamp 1571791925
transform 1 0 5842 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_402
timestamp 1571791925
transform 1 0 6670 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_403
timestamp 1571791925
transform 1 0 5934 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_404
timestamp 1571791925
transform 1 0 6854 0 1 8806
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_405
timestamp 1571791925
transform 1 0 6854 0 1 9486
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_406
timestamp 1571791925
transform 1 0 8970 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_407
timestamp 1571791925
transform 1 0 8970 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_408
timestamp 1571791925
transform 1 0 7958 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_409
timestamp 1571791925
transform 1 0 8602 0 1 8942
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_410
timestamp 1571791925
transform 1 0 8602 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_411
timestamp 1571791925
transform 1 0 8234 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_412
timestamp 1571791925
transform 1 0 9154 0 1 9554
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_413
timestamp 1571791925
transform 1 0 9246 0 1 8398
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_414
timestamp 1571791925
transform 1 0 8326 0 1 9486
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_415
timestamp 1571791925
transform 1 0 8510 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_416
timestamp 1571791925
transform 1 0 9430 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_417
timestamp 1571791925
transform 1 0 8878 0 1 8466
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_418
timestamp 1571791925
transform 1 0 8510 0 1 9350
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_419
timestamp 1571791925
transform 1 0 9246 0 1 10098
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_420
timestamp 1571791925
transform 1 0 9246 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_421
timestamp 1571791925
transform 1 0 8694 0 1 10234
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_422
timestamp 1571791925
transform 1 0 9338 0 1 9622
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_423
timestamp 1571791925
transform 1 0 9338 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_424
timestamp 1571791925
transform 1 0 8142 0 1 10506
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_425
timestamp 1571791925
transform 1 0 8418 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_426
timestamp 1571791925
transform 1 0 7866 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_427
timestamp 1571791925
transform 1 0 8510 0 1 10030
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_428
timestamp 1571791925
transform 1 0 8326 0 1 8874
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_429
timestamp 1571791925
transform 1 0 2346 0 1 5338
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_430
timestamp 1571791925
transform 1 0 5382 0 1 9962
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_431
timestamp 1571791925
transform 1 0 5382 0 1 4794
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_432
timestamp 1571791925
transform 1 0 2714 0 1 5338
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_433
timestamp 1571791925
transform 1 0 5382 0 1 7786
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_434
timestamp 1571791925
transform 1 0 2254 0 1 5338
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_435
timestamp 1571791925
transform 1 0 8234 0 1 12818
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_436
timestamp 1571791925
transform 1 0 7866 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_437
timestamp 1571791925
transform 1 0 9246 0 1 10982
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_438
timestamp 1571791925
transform 1 0 9338 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_439
timestamp 1571791925
transform 1 0 7866 0 1 11526
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_440
timestamp 1571791925
transform 1 0 9154 0 1 10982
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_441
timestamp 1571791925
transform 1 0 9338 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_442
timestamp 1571791925
transform 1 0 7958 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_443
timestamp 1571791925
transform 1 0 9154 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_444
timestamp 1571791925
transform 1 0 9246 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_445
timestamp 1571791925
transform 1 0 7958 0 1 12886
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_446
timestamp 1571791925
transform 1 0 8786 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_447
timestamp 1571791925
transform 1 0 8970 0 1 11050
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_448
timestamp 1571791925
transform 1 0 9430 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_449
timestamp 1571791925
transform 1 0 8602 0 1 12886
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_450
timestamp 1571791925
transform 1 0 9062 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_451
timestamp 1571791925
transform 1 0 9246 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_452
timestamp 1571791925
transform 1 0 8418 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_453
timestamp 1571791925
transform 1 0 8602 0 1 11322
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_454
timestamp 1571791925
transform 1 0 7774 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_455
timestamp 1571791925
transform 1 0 9338 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_456
timestamp 1571791925
transform 1 0 8326 0 1 12818
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_457
timestamp 1571791925
transform 1 0 6762 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_458
timestamp 1571791925
transform 1 0 6026 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_459
timestamp 1571791925
transform 1 0 6210 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_460
timestamp 1571791925
transform 1 0 5750 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_461
timestamp 1571791925
transform 1 0 5566 0 1 10982
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_462
timestamp 1571791925
transform 1 0 5934 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_463
timestamp 1571791925
transform 1 0 6854 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_464
timestamp 1571791925
transform 1 0 6394 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_465
timestamp 1571791925
transform 1 0 5934 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_466
timestamp 1571791925
transform 1 0 5842 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_467
timestamp 1571791925
transform 1 0 6394 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_468
timestamp 1571791925
transform 1 0 5566 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_469
timestamp 1571791925
transform 1 0 7130 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_470
timestamp 1571791925
transform 1 0 6486 0 1 12614
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_471
timestamp 1571791925
transform 1 0 5934 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_472
timestamp 1571791925
transform 1 0 7314 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_473
timestamp 1571791925
transform 1 0 6118 0 1 12954
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_474
timestamp 1571791925
transform 1 0 7406 0 1 14246
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_475
timestamp 1571791925
transform 1 0 7222 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_476
timestamp 1571791925
transform 1 0 5842 0 1 13974
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_477
timestamp 1571791925
transform 1 0 6854 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_478
timestamp 1571791925
transform 1 0 7038 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_479
timestamp 1571791925
transform 1 0 7222 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_480
timestamp 1571791925
transform 1 0 7038 0 1 14518
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_481
timestamp 1571791925
transform 1 0 7314 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_482
timestamp 1571791925
transform 1 0 6946 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_483
timestamp 1571791925
transform 1 0 7314 0 1 14246
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_484
timestamp 1571791925
transform 1 0 6670 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_485
timestamp 1571791925
transform 1 0 5842 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_486
timestamp 1571791925
transform 1 0 5842 0 1 15130
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_487
timestamp 1571791925
transform 1 0 6302 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_488
timestamp 1571791925
transform 1 0 5934 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_489
timestamp 1571791925
transform 1 0 5566 0 1 14042
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_490
timestamp 1571791925
transform 1 0 5934 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_491
timestamp 1571791925
transform 1 0 6578 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_492
timestamp 1571791925
transform 1 0 7222 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_493
timestamp 1571791925
transform 1 0 6486 0 1 15674
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_494
timestamp 1571791925
transform 1 0 6670 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_495
timestamp 1571791925
transform 1 0 6578 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_496
timestamp 1571791925
transform 1 0 7590 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_497
timestamp 1571791925
transform 1 0 8970 0 1 14790
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_498
timestamp 1571791925
transform 1 0 7682 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_499
timestamp 1571791925
transform 1 0 9246 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_500
timestamp 1571791925
transform 1 0 8786 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_501
timestamp 1571791925
transform 1 0 8510 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_502
timestamp 1571791925
transform 1 0 8418 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_503
timestamp 1571791925
transform 1 0 8602 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_504
timestamp 1571791925
transform 1 0 7590 0 1 13838
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_505
timestamp 1571791925
transform 1 0 9246 0 1 13974
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_506
timestamp 1571791925
transform 1 0 9246 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_507
timestamp 1571791925
transform 1 0 9154 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_508
timestamp 1571791925
transform 1 0 7774 0 1 15334
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_509
timestamp 1571791925
transform 1 0 8970 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_510
timestamp 1571791925
transform 1 0 9154 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_511
timestamp 1571791925
transform 1 0 7682 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_512
timestamp 1571791925
transform 1 0 4002 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_513
timestamp 1571791925
transform 1 0 4922 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_514
timestamp 1571791925
transform 1 0 5198 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_515
timestamp 1571791925
transform 1 0 4646 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_516
timestamp 1571791925
transform 1 0 4370 0 1 12818
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_517
timestamp 1571791925
transform 1 0 4646 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_518
timestamp 1571791925
transform 1 0 4738 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_519
timestamp 1571791925
transform 1 0 4922 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_520
timestamp 1571791925
transform 1 0 3818 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_521
timestamp 1571791925
transform 1 0 4554 0 1 11594
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_522
timestamp 1571791925
transform 1 0 3910 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_523
timestamp 1571791925
transform 1 0 5106 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_524
timestamp 1571791925
transform 1 0 4830 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_525
timestamp 1571791925
transform 1 0 4738 0 1 11798
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_526
timestamp 1571791925
transform 1 0 4094 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_527
timestamp 1571791925
transform 1 0 4646 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_528
timestamp 1571791925
transform 1 0 4186 0 1 12614
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_529
timestamp 1571791925
transform 1 0 5290 0 1 11526
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_530
timestamp 1571791925
transform 1 0 2898 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_531
timestamp 1571791925
transform 1 0 2438 0 1 12818
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_532
timestamp 1571791925
transform 1 0 1978 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_533
timestamp 1571791925
transform 1 0 2070 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_534
timestamp 1571791925
transform 1 0 1426 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_535
timestamp 1571791925
transform 1 0 1978 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_536
timestamp 1571791925
transform 1 0 2438 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_537
timestamp 1571791925
transform 1 0 2162 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_538
timestamp 1571791925
transform 1 0 2714 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_539
timestamp 1571791925
transform 1 0 2162 0 1 11526
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_540
timestamp 1571791925
transform 1 0 1702 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_541
timestamp 1571791925
transform 1 0 2070 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_542
timestamp 1571791925
transform 1 0 1518 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_543
timestamp 1571791925
transform 1 0 1794 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_544
timestamp 1571791925
transform 1 0 1702 0 1 11050
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_545
timestamp 1571791925
transform 1 0 3174 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_546
timestamp 1571791925
transform 1 0 3174 0 1 11322
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_547
timestamp 1571791925
transform 1 0 2346 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_548
timestamp 1571791925
transform 1 0 2806 0 1 11526
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_549
timestamp 1571791925
transform 1 0 2162 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_550
timestamp 1571791925
transform 1 0 1794 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_551
timestamp 1571791925
transform 1 0 2990 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_552
timestamp 1571791925
transform 1 0 1426 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_553
timestamp 1571791925
transform 1 0 1702 0 1 13362
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_554
timestamp 1571791925
transform 1 0 1794 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_555
timestamp 1571791925
transform 1 0 3174 0 1 13498
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_556
timestamp 1571791925
transform 1 0 2898 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_557
timestamp 1571791925
transform 1 0 1794 0 1 15538
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_558
timestamp 1571791925
transform 1 0 2162 0 1 14246
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_559
timestamp 1571791925
transform 1 0 2438 0 1 13838
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_560
timestamp 1571791925
transform 1 0 2346 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_561
timestamp 1571791925
transform 1 0 3174 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_562
timestamp 1571791925
transform 1 0 2346 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_563
timestamp 1571791925
transform 1 0 2806 0 1 14858
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_564
timestamp 1571791925
transform 1 0 1978 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_565
timestamp 1571791925
transform 1 0 2898 0 1 13974
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_566
timestamp 1571791925
transform 1 0 2070 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_567
timestamp 1571791925
transform 1 0 1518 0 1 15130
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_568
timestamp 1571791925
transform 1 0 2714 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_569
timestamp 1571791925
transform 1 0 2070 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_570
timestamp 1571791925
transform 1 0 2070 0 1 14246
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_571
timestamp 1571791925
transform 1 0 2346 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_572
timestamp 1571791925
transform 1 0 4462 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_573
timestamp 1571791925
transform 1 0 4830 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_574
timestamp 1571791925
transform 1 0 4186 0 1 15538
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_575
timestamp 1571791925
transform 1 0 3450 0 1 15130
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_576
timestamp 1571791925
transform 1 0 4186 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_577
timestamp 1571791925
transform 1 0 4554 0 1 13362
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_578
timestamp 1571791925
transform 1 0 4738 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_579
timestamp 1571791925
transform 1 0 5014 0 1 15538
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_580
timestamp 1571791925
transform 1 0 3542 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_581
timestamp 1571791925
transform 1 0 4462 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_582
timestamp 1571791925
transform 1 0 5198 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_583
timestamp 1571791925
transform 1 0 3542 0 1 15674
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_584
timestamp 1571791925
transform 1 0 3726 0 1 13838
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_585
timestamp 1571791925
transform 1 0 5198 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_586
timestamp 1571791925
transform 1 0 3542 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_587
timestamp 1571791925
transform 1 0 3358 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_588
timestamp 1571791925
transform 1 0 5198 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_589
timestamp 1571791925
transform 1 0 3634 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_590
timestamp 1571791925
transform 1 0 4554 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_591
timestamp 1571791925
transform 1 0 5106 0 1 18326
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_592
timestamp 1571791925
transform 1 0 4186 0 1 16422
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_593
timestamp 1571791925
transform 1 0 3818 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_594
timestamp 1571791925
transform 1 0 5106 0 1 17714
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_595
timestamp 1571791925
transform 1 0 4738 0 1 16490
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_596
timestamp 1571791925
transform 1 0 3818 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_597
timestamp 1571791925
transform 1 0 3450 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_598
timestamp 1571791925
transform 1 0 4646 0 1 16014
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_599
timestamp 1571791925
transform 1 0 4830 0 1 17646
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_600
timestamp 1571791925
transform 1 0 3726 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_601
timestamp 1571791925
transform 1 0 4830 0 1 18394
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_602
timestamp 1571791925
transform 1 0 4370 0 1 16014
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_603
timestamp 1571791925
transform 1 0 4002 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_604
timestamp 1571791925
transform 1 0 4186 0 1 16014
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_605
timestamp 1571791925
transform 1 0 4002 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_606
timestamp 1571791925
transform 1 0 4370 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_607
timestamp 1571791925
transform 1 0 3818 0 1 17714
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_608
timestamp 1571791925
transform 1 0 3082 0 1 16150
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_609
timestamp 1571791925
transform 1 0 1518 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_610
timestamp 1571791925
transform 1 0 1518 0 1 17850
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_611
timestamp 1571791925
transform 1 0 2162 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_612
timestamp 1571791925
transform 1 0 3266 0 1 17714
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_613
timestamp 1571791925
transform 1 0 3082 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_614
timestamp 1571791925
transform 1 0 1426 0 1 16626
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_615
timestamp 1571791925
transform 1 0 1610 0 1 18054
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_616
timestamp 1571791925
transform 1 0 2990 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_617
timestamp 1571791925
transform 1 0 2898 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_618
timestamp 1571791925
transform 1 0 2714 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_619
timestamp 1571791925
transform 1 0 1702 0 1 16490
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_620
timestamp 1571791925
transform 1 0 3174 0 1 16422
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_621
timestamp 1571791925
transform 1 0 2070 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_622
timestamp 1571791925
transform 1 0 2530 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_623
timestamp 1571791925
transform 1 0 2898 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_624
timestamp 1571791925
transform 1 0 2806 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_625
timestamp 1571791925
transform 1 0 2530 0 1 16150
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_626
timestamp 1571791925
transform 1 0 3266 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_627
timestamp 1571791925
transform 1 0 2070 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_628
timestamp 1571791925
transform 1 0 2162 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_629
timestamp 1571791925
transform 1 0 2254 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_630
timestamp 1571791925
transform 1 0 1978 0 1 18666
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_631
timestamp 1571791925
transform 1 0 4554 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_632
timestamp 1571791925
transform 1 0 4370 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_633
timestamp 1571791925
transform 1 0 4186 0 1 18598
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_634
timestamp 1571791925
transform 1 0 3358 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_635
timestamp 1571791925
transform 1 0 6762 0 1 17102
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_636
timestamp 1571791925
transform 1 0 9154 0 1 16626
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_637
timestamp 1571791925
transform 1 0 9430 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_638
timestamp 1571791925
transform 1 0 9062 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_639
timestamp 1571791925
transform 1 0 9062 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_640
timestamp 1571791925
transform 1 0 9338 0 1 16966
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_641
timestamp 1571791925
transform 1 0 8786 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_642
timestamp 1571791925
transform 1 0 9154 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_643
timestamp 1571791925
transform 1 0 8878 0 1 16014
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_644
timestamp 1571791925
transform 1 0 6210 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_645
timestamp 1571791925
transform 1 0 6486 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_646
timestamp 1571791925
transform 1 0 5750 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_647
timestamp 1571791925
transform 1 0 6118 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_648
timestamp 1571791925
transform 1 0 7038 0 1 17102
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_649
timestamp 1571791925
transform 1 0 6026 0 1 16626
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_650
timestamp 1571791925
transform 1 0 5842 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_651
timestamp 1571791925
transform 1 0 8970 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_652
timestamp 1571791925
transform 1 0 9338 0 1 17510
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_653
timestamp 1571791925
transform 1 0 9430 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_654
timestamp 1571791925
transform 1 0 5566 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_655
timestamp 1571791925
transform 1 0 8970 0 1 17782
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_656
timestamp 1571791925
transform 1 0 8786 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_657
timestamp 1571791925
transform 1 0 7682 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_658
timestamp 1571791925
transform 1 0 5658 0 1 18122
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_659
timestamp 1571791925
transform 1 0 6026 0 1 18394
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_660
timestamp 1571791925
transform 1 0 8326 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_661
timestamp 1571791925
transform 1 0 8234 0 1 18598
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_662
timestamp 1571791925
transform 1 0 6486 0 1 18054
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_663
timestamp 1571791925
transform 1 0 7774 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_664
timestamp 1571791925
transform 1 0 6118 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_665
timestamp 1571791925
transform 1 0 6854 0 1 17510
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_666
timestamp 1571791925
transform 1 0 6670 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_667
timestamp 1571791925
transform 1 0 6762 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_668
timestamp 1571791925
transform 1 0 6118 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_669
timestamp 1571791925
transform 1 0 5934 0 1 18394
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_670
timestamp 1571791925
transform 1 0 9246 0 1 17510
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_671
timestamp 1571791925
transform 1 0 9246 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_672
timestamp 1571791925
transform 1 0 6578 0 1 18258
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_673
timestamp 1571791925
transform 1 0 9430 0 1 16490
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_674
timestamp 1571791925
transform 1 0 7774 0 1 17646
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_675
timestamp 1571791925
transform 1 0 7314 0 1 18054
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_676
timestamp 1571791925
transform 1 0 8694 0 1 17102
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_677
timestamp 1571791925
transform 1 0 8510 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_678
timestamp 1571791925
transform 1 0 8878 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_679
timestamp 1571791925
transform 1 0 6946 0 1 16626
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_680
timestamp 1571791925
transform 1 0 5382 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_681
timestamp 1571791925
transform 1 0 5382 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_682
timestamp 1571791925
transform 1 0 5382 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_683
timestamp 1571791925
transform 1 0 5382 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_684
timestamp 1571791925
transform 1 0 16882 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_685
timestamp 1571791925
transform 1 0 16698 0 1 11594
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_686
timestamp 1571791925
transform 1 0 17066 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_687
timestamp 1571791925
transform 1 0 17250 0 1 11798
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_688
timestamp 1571791925
transform 1 0 17710 0 1 11798
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_689
timestamp 1571791925
transform 1 0 17526 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_690
timestamp 1571791925
transform 1 0 16422 0 1 12614
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_691
timestamp 1571791925
transform 1 0 16238 0 1 11254
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_692
timestamp 1571791925
transform 1 0 17434 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_693
timestamp 1571791925
transform 1 0 17250 0 1 11050
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_694
timestamp 1571791925
transform 1 0 17342 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_695
timestamp 1571791925
transform 1 0 16698 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_696
timestamp 1571791925
transform 1 0 16974 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_697
timestamp 1571791925
transform 1 0 15318 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_698
timestamp 1571791925
transform 1 0 14490 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_699
timestamp 1571791925
transform 1 0 15410 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_700
timestamp 1571791925
transform 1 0 15134 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_701
timestamp 1571791925
transform 1 0 14766 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_702
timestamp 1571791925
transform 1 0 14950 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_703
timestamp 1571791925
transform 1 0 14214 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_704
timestamp 1571791925
transform 1 0 15410 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_705
timestamp 1571791925
transform 1 0 15502 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_706
timestamp 1571791925
transform 1 0 15042 0 1 11798
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_707
timestamp 1571791925
transform 1 0 14674 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_708
timestamp 1571791925
transform 1 0 14766 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_709
timestamp 1571791925
transform 1 0 13754 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_710
timestamp 1571791925
transform 1 0 14766 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_711
timestamp 1571791925
transform 1 0 13938 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_712
timestamp 1571791925
transform 1 0 13754 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_713
timestamp 1571791925
transform 1 0 14122 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_714
timestamp 1571791925
transform 1 0 15134 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_715
timestamp 1571791925
transform 1 0 15318 0 1 15130
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_716
timestamp 1571791925
transform 1 0 15594 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_717
timestamp 1571791925
transform 1 0 15594 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_718
timestamp 1571791925
transform 1 0 14306 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_719
timestamp 1571791925
transform 1 0 14674 0 1 14790
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_720
timestamp 1571791925
transform 1 0 15226 0 1 15130
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_721
timestamp 1571791925
transform 1 0 15410 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_722
timestamp 1571791925
transform 1 0 15502 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_723
timestamp 1571791925
transform 1 0 15318 0 1 13430
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_724
timestamp 1571791925
transform 1 0 15134 0 1 13974
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_725
timestamp 1571791925
transform 1 0 15134 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_726
timestamp 1571791925
transform 1 0 14214 0 1 15334
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_727
timestamp 1571791925
transform 1 0 14398 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_728
timestamp 1571791925
transform 1 0 14950 0 1 14858
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_729
timestamp 1571791925
transform 1 0 16422 0 1 14586
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_730
timestamp 1571791925
transform 1 0 16054 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_731
timestamp 1571791925
transform 1 0 15870 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_732
timestamp 1571791925
transform 1 0 15870 0 1 14246
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_733
timestamp 1571791925
transform 1 0 16238 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_734
timestamp 1571791925
transform 1 0 15686 0 1 13158
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_735
timestamp 1571791925
transform 1 0 15686 0 1 14790
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_736
timestamp 1571791925
transform 1 0 13386 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_737
timestamp 1571791925
transform 1 0 13294 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_738
timestamp 1571791925
transform 1 0 11822 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_739
timestamp 1571791925
transform 1 0 12098 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_740
timestamp 1571791925
transform 1 0 13018 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_741
timestamp 1571791925
transform 1 0 13570 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_742
timestamp 1571791925
transform 1 0 13202 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_743
timestamp 1571791925
transform 1 0 12190 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_744
timestamp 1571791925
transform 1 0 13386 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_745
timestamp 1571791925
transform 1 0 12650 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_746
timestamp 1571791925
transform 1 0 12558 0 1 11730
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_747
timestamp 1571791925
transform 1 0 12098 0 1 12138
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_748
timestamp 1571791925
transform 1 0 12466 0 1 12342
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_749
timestamp 1571791925
transform 1 0 13294 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_750
timestamp 1571791925
transform 1 0 12834 0 1 12070
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_751
timestamp 1571791925
transform 1 0 12282 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_752
timestamp 1571791925
transform 1 0 12742 0 1 12070
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_753
timestamp 1571791925
transform 1 0 13570 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_754
timestamp 1571791925
transform 1 0 12558 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_755
timestamp 1571791925
transform 1 0 12190 0 1 11050
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_756
timestamp 1571791925
transform 1 0 12926 0 1 10710
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_757
timestamp 1571791925
transform 1 0 12926 0 1 11118
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_758
timestamp 1571791925
transform 1 0 13018 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_759
timestamp 1571791925
transform 1 0 12374 0 1 12274
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_760
timestamp 1571791925
transform 1 0 13386 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_761
timestamp 1571791925
transform 1 0 13294 0 1 11662
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_762
timestamp 1571791925
transform 1 0 10810 0 1 10778
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_763
timestamp 1571791925
transform 1 0 10718 0 1 10642
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_764
timestamp 1571791925
transform 1 0 10074 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_765
timestamp 1571791925
transform 1 0 9798 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_766
timestamp 1571791925
transform 1 0 10258 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_767
timestamp 1571791925
transform 1 0 11086 0 1 12750
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_768
timestamp 1571791925
transform 1 0 10074 0 1 12682
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_769
timestamp 1571791925
transform 1 0 11362 0 1 13226
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_770
timestamp 1571791925
transform 1 0 10626 0 1 12410
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_771
timestamp 1571791925
transform 1 0 9982 0 1 11050
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_772
timestamp 1571791925
transform 1 0 11454 0 1 10982
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_773
timestamp 1571791925
transform 1 0 9982 0 1 12206
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_774
timestamp 1571791925
transform 1 0 9706 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_775
timestamp 1571791925
transform 1 0 10994 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_776
timestamp 1571791925
transform 1 0 10258 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_777
timestamp 1571791925
transform 1 0 11086 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_778
timestamp 1571791925
transform 1 0 11270 0 1 14790
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_779
timestamp 1571791925
transform 1 0 10258 0 1 15334
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_780
timestamp 1571791925
transform 1 0 10350 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_781
timestamp 1571791925
transform 1 0 11178 0 1 14994
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_782
timestamp 1571791925
transform 1 0 10534 0 1 14314
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_783
timestamp 1571791925
transform 1 0 11178 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_784
timestamp 1571791925
transform 1 0 11454 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_785
timestamp 1571791925
transform 1 0 10718 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_786
timestamp 1571791925
transform 1 0 10074 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_787
timestamp 1571791925
transform 1 0 11638 0 1 13838
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_788
timestamp 1571791925
transform 1 0 11730 0 1 15062
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_789
timestamp 1571791925
transform 1 0 12190 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_790
timestamp 1571791925
transform 1 0 12742 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_791
timestamp 1571791925
transform 1 0 11730 0 1 15334
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_792
timestamp 1571791925
transform 1 0 11638 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_793
timestamp 1571791925
transform 1 0 13294 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_794
timestamp 1571791925
transform 1 0 11730 0 1 13906
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_795
timestamp 1571791925
transform 1 0 12558 0 1 15470
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_796
timestamp 1571791925
transform 1 0 12282 0 1 14586
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_797
timestamp 1571791925
transform 1 0 11840 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_798
timestamp 1571791925
transform 1 0 12006 0 1 15402
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_799
timestamp 1571791925
transform 1 0 13018 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_800
timestamp 1571791925
transform 1 0 12650 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_801
timestamp 1571791925
transform 1 0 12558 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_802
timestamp 1571791925
transform 1 0 12006 0 1 14450
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_803
timestamp 1571791925
transform 1 0 12466 0 1 14382
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_804
timestamp 1571791925
transform 1 0 12834 0 1 14586
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_805
timestamp 1571791925
transform 1 0 13202 0 1 15062
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_806
timestamp 1571791925
transform 1 0 13202 0 1 15334
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_807
timestamp 1571791925
transform 1 0 12006 0 1 13362
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_808
timestamp 1571791925
transform 1 0 13202 0 1 13702
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_809
timestamp 1571791925
transform 1 0 12926 0 1 14926
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_810
timestamp 1571791925
transform 1 0 11546 0 1 12886
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_811
timestamp 1571791925
transform 1 0 11546 0 1 11866
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_812
timestamp 1571791925
transform 1 0 11546 0 1 13294
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_813
timestamp 1571791925
transform 1 0 11546 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_814
timestamp 1571791925
transform 1 0 12190 0 1 17646
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_815
timestamp 1571791925
transform 1 0 10902 0 1 16762
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_816
timestamp 1571791925
transform 1 0 9614 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_817
timestamp 1571791925
transform 1 0 13294 0 1 16966
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_818
timestamp 1571791925
transform 1 0 11822 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_819
timestamp 1571791925
transform 1 0 11914 0 1 17510
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_820
timestamp 1571791925
transform 1 0 11178 0 1 18054
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_821
timestamp 1571791925
transform 1 0 12006 0 1 17714
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_822
timestamp 1571791925
transform 1 0 10442 0 1 17714
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_823
timestamp 1571791925
transform 1 0 10902 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_824
timestamp 1571791925
transform 1 0 11546 0 1 17102
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_825
timestamp 1571791925
transform 1 0 10902 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_826
timestamp 1571791925
transform 1 0 12374 0 1 17510
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_827
timestamp 1571791925
transform 1 0 11362 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_828
timestamp 1571791925
transform 1 0 11270 0 1 17646
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_829
timestamp 1571791925
transform 1 0 10534 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_830
timestamp 1571791925
transform 1 0 10902 0 1 17646
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_831
timestamp 1571791925
transform 1 0 9890 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_832
timestamp 1571791925
transform 1 0 10350 0 1 17238
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_833
timestamp 1571791925
transform 1 0 9706 0 1 18190
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_834
timestamp 1571791925
transform 1 0 10534 0 1 18598
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_835
timestamp 1571791925
transform 1 0 12650 0 1 16762
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_836
timestamp 1571791925
transform 1 0 10258 0 1 16218
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_837
timestamp 1571791925
transform 1 0 10994 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_838
timestamp 1571791925
transform 1 0 10626 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_839
timestamp 1571791925
transform 1 0 12558 0 1 16558
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_840
timestamp 1571791925
transform 1 0 10166 0 1 16082
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_841
timestamp 1571791925
transform 1 0 10442 0 1 18734
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_842
timestamp 1571791925
transform 1 0 11178 0 1 17170
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_843
timestamp 1571791925
transform 1 0 10718 0 1 17306
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_844
timestamp 1571791925
transform 1 0 12834 0 1 15878
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_845
timestamp 1571791925
transform 1 0 9522 0 1 3026
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_846
timestamp 1571791925
transform 1 0 9522 0 1 17578
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_847
timestamp 1571791925
transform 1 0 9522 0 1 11186
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_848
timestamp 1571791925
transform 1 0 9522 0 1 3366
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_849
timestamp 1571791925
transform 1 0 9522 0 1 8602
box -29 -23 29 23
use VIA_L1M1_PR_MR  VIA_L1M1_PR_MR_850
timestamp 1571791925
transform 1 0 9522 0 1 13226
box -29 -23 29 23
use VIA_M1M2_PR  VIA_M1M2_PR_0
timestamp 1571791925
transform 1 0 13754 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_1
timestamp 1571791925
transform 1 0 15778 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_2
timestamp 1571791925
transform 1 0 13754 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_3
timestamp 1571791925
transform 1 0 15778 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_4
timestamp 1571791925
transform 1 0 14950 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_5
timestamp 1571791925
transform 1 0 14950 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_6
timestamp 1571791925
transform 1 0 15502 0 1 2958
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_7
timestamp 1571791925
transform 1 0 13662 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_8
timestamp 1571791925
transform 1 0 14306 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_9
timestamp 1571791925
transform 1 0 14398 0 1 2550
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_10
timestamp 1571791925
transform 1 0 14398 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_11
timestamp 1571791925
transform 1 0 15502 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_12
timestamp 1571791925
transform 1 0 15410 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_13
timestamp 1571791925
transform 1 0 15410 0 1 4522
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_14
timestamp 1571791925
transform 1 0 13938 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_15
timestamp 1571791925
transform 1 0 13938 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_16
timestamp 1571791925
transform 1 0 14398 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_17
timestamp 1571791925
transform 1 0 14858 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_18
timestamp 1571791925
transform 1 0 13754 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_19
timestamp 1571791925
transform 1 0 15042 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_20
timestamp 1571791925
transform 1 0 13662 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_21
timestamp 1571791925
transform 1 0 14858 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_22
timestamp 1571791925
transform 1 0 14858 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_23
timestamp 1571791925
transform 1 0 15962 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_24
timestamp 1571791925
transform 1 0 15962 0 1 3162
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_25
timestamp 1571791925
transform 1 0 13754 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_26
timestamp 1571791925
transform 1 0 13662 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_27
timestamp 1571791925
transform 1 0 13662 0 1 3162
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_28
timestamp 1571791925
transform 1 0 14306 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_29
timestamp 1571791925
transform 1 0 13846 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_30
timestamp 1571791925
transform 1 0 13846 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_31
timestamp 1571791925
transform 1 0 15778 0 1 4454
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_32
timestamp 1571791925
transform 1 0 14306 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_33
timestamp 1571791925
transform 1 0 12374 0 1 2618
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_34
timestamp 1571791925
transform 1 0 12466 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_35
timestamp 1571791925
transform 1 0 12926 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_36
timestamp 1571791925
transform 1 0 9982 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_37
timestamp 1571791925
transform 1 0 9706 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_38
timestamp 1571791925
transform 1 0 11454 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_39
timestamp 1571791925
transform 1 0 10902 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_40
timestamp 1571791925
transform 1 0 10626 0 1 3910
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_41
timestamp 1571791925
transform 1 0 10534 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_42
timestamp 1571791925
transform 1 0 10718 0 1 4794
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_43
timestamp 1571791925
transform 1 0 9614 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_44
timestamp 1571791925
transform 1 0 10626 0 1 5066
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_45
timestamp 1571791925
transform 1 0 10626 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_46
timestamp 1571791925
transform 1 0 9614 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_47
timestamp 1571791925
transform 1 0 10810 0 1 3162
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_48
timestamp 1571791925
transform 1 0 9614 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_49
timestamp 1571791925
transform 1 0 9982 0 1 3706
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_50
timestamp 1571791925
transform 1 0 10534 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_51
timestamp 1571791925
transform 1 0 11454 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_52
timestamp 1571791925
transform 1 0 9982 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_53
timestamp 1571791925
transform 1 0 9798 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_54
timestamp 1571791925
transform 1 0 10258 0 1 3638
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_55
timestamp 1571791925
transform 1 0 10258 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_56
timestamp 1571791925
transform 1 0 9798 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_57
timestamp 1571791925
transform 1 0 10902 0 1 4658
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_58
timestamp 1571791925
transform 1 0 9706 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_59
timestamp 1571791925
transform 1 0 13294 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_60
timestamp 1571791925
transform 1 0 13294 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_61
timestamp 1571791925
transform 1 0 12926 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_62
timestamp 1571791925
transform 1 0 12374 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_63
timestamp 1571791925
transform 1 0 11638 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_64
timestamp 1571791925
transform 1 0 13386 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_65
timestamp 1571791925
transform 1 0 13386 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_66
timestamp 1571791925
transform 1 0 12834 0 1 4046
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_67
timestamp 1571791925
transform 1 0 11638 0 1 4658
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_68
timestamp 1571791925
transform 1 0 11730 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_69
timestamp 1571791925
transform 1 0 12282 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_70
timestamp 1571791925
transform 1 0 11638 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_71
timestamp 1571791925
transform 1 0 11730 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_72
timestamp 1571791925
transform 1 0 13570 0 1 4046
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_73
timestamp 1571791925
transform 1 0 13478 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_74
timestamp 1571791925
transform 1 0 11914 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_75
timestamp 1571791925
transform 1 0 11914 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_76
timestamp 1571791925
transform 1 0 11546 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_77
timestamp 1571791925
transform 1 0 13478 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_78
timestamp 1571791925
transform 1 0 12558 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_79
timestamp 1571791925
transform 1 0 13018 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_80
timestamp 1571791925
transform 1 0 13018 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_81
timestamp 1571791925
transform 1 0 11822 0 1 6902
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_82
timestamp 1571791925
transform 1 0 11822 0 1 7310
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_83
timestamp 1571791925
transform 1 0 12282 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_84
timestamp 1571791925
transform 1 0 13294 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_85
timestamp 1571791925
transform 1 0 13294 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_86
timestamp 1571791925
transform 1 0 12650 0 1 6086
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_87
timestamp 1571791925
transform 1 0 12650 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_88
timestamp 1571791925
transform 1 0 12834 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_89
timestamp 1571791925
transform 1 0 12282 0 1 7718
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_90
timestamp 1571791925
transform 1 0 12282 0 1 7446
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_91
timestamp 1571791925
transform 1 0 13018 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_92
timestamp 1571791925
transform 1 0 13110 0 1 5814
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_93
timestamp 1571791925
transform 1 0 13110 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_94
timestamp 1571791925
transform 1 0 11638 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_95
timestamp 1571791925
transform 1 0 12558 0 1 7718
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_96
timestamp 1571791925
transform 1 0 12098 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_97
timestamp 1571791925
transform 1 0 13570 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_98
timestamp 1571791925
transform 1 0 13294 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_99
timestamp 1571791925
transform 1 0 12098 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_100
timestamp 1571791925
transform 1 0 10810 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_101
timestamp 1571791925
transform 1 0 11362 0 1 5746
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_102
timestamp 1571791925
transform 1 0 11178 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_103
timestamp 1571791925
transform 1 0 11362 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_104
timestamp 1571791925
transform 1 0 10350 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_105
timestamp 1571791925
transform 1 0 10350 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_106
timestamp 1571791925
transform 1 0 10902 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_107
timestamp 1571791925
transform 1 0 11362 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_108
timestamp 1571791925
transform 1 0 10902 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_109
timestamp 1571791925
transform 1 0 11454 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_110
timestamp 1571791925
transform 1 0 11270 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_111
timestamp 1571791925
transform 1 0 10626 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_112
timestamp 1571791925
transform 1 0 10626 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_113
timestamp 1571791925
transform 1 0 11270 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_114
timestamp 1571791925
transform 1 0 10718 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_115
timestamp 1571791925
transform 1 0 11178 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_116
timestamp 1571791925
transform 1 0 10074 0 1 5746
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_117
timestamp 1571791925
transform 1 0 10534 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_118
timestamp 1571791925
transform 1 0 11454 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_119
timestamp 1571791925
transform 1 0 11454 0 1 6630
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_120
timestamp 1571791925
transform 1 0 10074 0 1 6154
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_121
timestamp 1571791925
transform 1 0 10718 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_122
timestamp 1571791925
transform 1 0 9890 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_123
timestamp 1571791925
transform 1 0 10718 0 1 6834
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_124
timestamp 1571791925
transform 1 0 9982 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_125
timestamp 1571791925
transform 1 0 9614 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_126
timestamp 1571791925
transform 1 0 11454 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_127
timestamp 1571791925
transform 1 0 10074 0 1 9350
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_128
timestamp 1571791925
transform 1 0 10810 0 1 9146
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_129
timestamp 1571791925
transform 1 0 10074 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_130
timestamp 1571791925
transform 1 0 11454 0 1 9010
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_131
timestamp 1571791925
transform 1 0 10718 0 1 9146
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_132
timestamp 1571791925
transform 1 0 10718 0 1 9486
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_133
timestamp 1571791925
transform 1 0 10718 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_134
timestamp 1571791925
transform 1 0 9982 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_135
timestamp 1571791925
transform 1 0 10626 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_136
timestamp 1571791925
transform 1 0 9890 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_137
timestamp 1571791925
transform 1 0 10626 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_138
timestamp 1571791925
transform 1 0 11362 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_139
timestamp 1571791925
transform 1 0 9982 0 1 9350
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_140
timestamp 1571791925
transform 1 0 9614 0 1 9010
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_141
timestamp 1571791925
transform 1 0 10994 0 1 10506
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_142
timestamp 1571791925
transform 1 0 10994 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_143
timestamp 1571791925
transform 1 0 11730 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_144
timestamp 1571791925
transform 1 0 12466 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_145
timestamp 1571791925
transform 1 0 11730 0 1 9962
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_146
timestamp 1571791925
transform 1 0 12098 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_147
timestamp 1571791925
transform 1 0 12466 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_148
timestamp 1571791925
transform 1 0 12834 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_149
timestamp 1571791925
transform 1 0 13018 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_150
timestamp 1571791925
transform 1 0 12834 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_151
timestamp 1571791925
transform 1 0 12006 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_152
timestamp 1571791925
transform 1 0 12558 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_153
timestamp 1571791925
transform 1 0 11546 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_154
timestamp 1571791925
transform 1 0 11546 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_155
timestamp 1571791925
transform 1 0 16790 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_156
timestamp 1571791925
transform 1 0 17434 0 1 7922
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_157
timestamp 1571791925
transform 1 0 17618 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_158
timestamp 1571791925
transform 1 0 14398 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_159
timestamp 1571791925
transform 1 0 14398 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_160
timestamp 1571791925
transform 1 0 14214 0 1 6630
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_161
timestamp 1571791925
transform 1 0 14214 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_162
timestamp 1571791925
transform 1 0 14398 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_163
timestamp 1571791925
transform 1 0 14306 0 1 7718
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_164
timestamp 1571791925
transform 1 0 14306 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_165
timestamp 1571791925
transform 1 0 13846 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_166
timestamp 1571791925
transform 1 0 13662 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_167
timestamp 1571791925
transform 1 0 13662 0 1 6630
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_168
timestamp 1571791925
transform 1 0 15042 0 1 6086
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_169
timestamp 1571791925
transform 1 0 15042 0 1 5746
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_170
timestamp 1571791925
transform 1 0 14490 0 1 7922
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_171
timestamp 1571791925
transform 1 0 15410 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_172
timestamp 1571791925
transform 1 0 14398 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_173
timestamp 1571791925
transform 1 0 15410 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_174
timestamp 1571791925
transform 1 0 15502 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_175
timestamp 1571791925
transform 1 0 15502 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_176
timestamp 1571791925
transform 1 0 15594 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_177
timestamp 1571791925
transform 1 0 15594 0 1 9962
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_178
timestamp 1571791925
transform 1 0 14490 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_179
timestamp 1571791925
transform 1 0 15410 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_180
timestamp 1571791925
transform 1 0 15410 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_181
timestamp 1571791925
transform 1 0 14490 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_182
timestamp 1571791925
transform 1 0 14490 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_183
timestamp 1571791925
transform 1 0 14766 0 1 9010
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_184
timestamp 1571791925
transform 1 0 14766 0 1 9418
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_185
timestamp 1571791925
transform 1 0 14950 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_186
timestamp 1571791925
transform 1 0 14950 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_187
timestamp 1571791925
transform 1 0 17158 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_188
timestamp 1571791925
transform 1 0 16790 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_189
timestamp 1571791925
transform 1 0 17526 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_190
timestamp 1571791925
transform 1 0 17618 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_191
timestamp 1571791925
transform 1 0 17342 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_192
timestamp 1571791925
transform 1 0 17434 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_193
timestamp 1571791925
transform 1 0 17526 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_194
timestamp 1571791925
transform 1 0 17526 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_195
timestamp 1571791925
transform 1 0 17434 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_196
timestamp 1571791925
transform 1 0 16698 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_197
timestamp 1571791925
transform 1 0 16698 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_198
timestamp 1571791925
transform 1 0 17526 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_199
timestamp 1571791925
transform 1 0 16146 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_200
timestamp 1571791925
transform 1 0 16146 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_201
timestamp 1571791925
transform 1 0 16698 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_202
timestamp 1571791925
transform 1 0 16698 0 1 9690
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_203
timestamp 1571791925
transform 1 0 16514 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_204
timestamp 1571791925
transform 1 0 16514 0 1 9894
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_205
timestamp 1571791925
transform 1 0 15686 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_206
timestamp 1571791925
transform 1 0 15686 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_207
timestamp 1571791925
transform 1 0 12834 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_208
timestamp 1571791925
transform 1 0 13846 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_209
timestamp 1571791925
transform 1 0 7682 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_210
timestamp 1571791925
transform 1 0 8234 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_211
timestamp 1571791925
transform 1 0 9154 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_212
timestamp 1571791925
transform 1 0 7590 0 1 2618
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_213
timestamp 1571791925
transform 1 0 7222 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_214
timestamp 1571791925
transform 1 0 6394 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_215
timestamp 1571791925
transform 1 0 6762 0 1 2482
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_216
timestamp 1571791925
transform 1 0 7130 0 1 2618
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_217
timestamp 1571791925
transform 1 0 6670 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_218
timestamp 1571791925
transform 1 0 6210 0 1 3162
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_219
timestamp 1571791925
transform 1 0 7406 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_220
timestamp 1571791925
transform 1 0 6210 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_221
timestamp 1571791925
transform 1 0 5842 0 1 5066
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_222
timestamp 1571791925
transform 1 0 6302 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_223
timestamp 1571791925
transform 1 0 7222 0 1 2958
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_224
timestamp 1571791925
transform 1 0 6302 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_225
timestamp 1571791925
transform 1 0 5750 0 1 2958
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_226
timestamp 1571791925
transform 1 0 5474 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_227
timestamp 1571791925
transform 1 0 6210 0 1 4794
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_228
timestamp 1571791925
transform 1 0 5658 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_229
timestamp 1571791925
transform 1 0 7130 0 1 3434
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_230
timestamp 1571791925
transform 1 0 5474 0 1 3706
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_231
timestamp 1571791925
transform 1 0 6854 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_232
timestamp 1571791925
transform 1 0 5842 0 1 4658
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_233
timestamp 1571791925
transform 1 0 5658 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_234
timestamp 1571791925
transform 1 0 5566 0 1 4794
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_235
timestamp 1571791925
transform 1 0 6762 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_236
timestamp 1571791925
transform 1 0 6670 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_237
timestamp 1571791925
transform 1 0 6486 0 1 3978
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_238
timestamp 1571791925
transform 1 0 6946 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_239
timestamp 1571791925
transform 1 0 6946 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_240
timestamp 1571791925
transform 1 0 6210 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_241
timestamp 1571791925
transform 1 0 6486 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_242
timestamp 1571791925
transform 1 0 5750 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_243
timestamp 1571791925
transform 1 0 6394 0 1 4250
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_244
timestamp 1571791925
transform 1 0 7682 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_245
timestamp 1571791925
transform 1 0 7590 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_246
timestamp 1571791925
transform 1 0 7866 0 1 4522
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_247
timestamp 1571791925
transform 1 0 7498 0 1 4522
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_248
timestamp 1571791925
transform 1 0 7866 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_249
timestamp 1571791925
transform 1 0 8510 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_250
timestamp 1571791925
transform 1 0 8970 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_251
timestamp 1571791925
transform 1 0 7774 0 1 4250
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_252
timestamp 1571791925
transform 1 0 9246 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_253
timestamp 1571791925
transform 1 0 9246 0 1 4794
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_254
timestamp 1571791925
transform 1 0 9154 0 1 2958
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_255
timestamp 1571791925
transform 1 0 7682 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_256
timestamp 1571791925
transform 1 0 7682 0 1 3162
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_257
timestamp 1571791925
transform 1 0 8050 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_258
timestamp 1571791925
transform 1 0 7774 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_259
timestamp 1571791925
transform 1 0 8694 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_260
timestamp 1571791925
transform 1 0 8234 0 1 4658
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_261
timestamp 1571791925
transform 1 0 8694 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_262
timestamp 1571791925
transform 1 0 8234 0 1 4046
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_263
timestamp 1571791925
transform 1 0 8234 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_264
timestamp 1571791925
transform 1 0 8234 0 1 3706
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_265
timestamp 1571791925
transform 1 0 3450 0 1 2618
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_266
timestamp 1571791925
transform 1 0 3542 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_267
timestamp 1571791925
transform 1 0 2530 0 1 2618
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_268
timestamp 1571791925
transform 1 0 2162 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_269
timestamp 1571791925
transform 1 0 1978 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_270
timestamp 1571791925
transform 1 0 2622 0 1 2414
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_271
timestamp 1571791925
transform 1 0 1426 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_272
timestamp 1571791925
transform 1 0 1978 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_273
timestamp 1571791925
transform 1 0 2990 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_274
timestamp 1571791925
transform 1 0 1794 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_275
timestamp 1571791925
transform 1 0 2346 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_276
timestamp 1571791925
transform 1 0 2346 0 1 3910
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_277
timestamp 1571791925
transform 1 0 1978 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_278
timestamp 1571791925
transform 1 0 1978 0 1 3366
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_279
timestamp 1571791925
transform 1 0 1702 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_280
timestamp 1571791925
transform 1 0 1794 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_281
timestamp 1571791925
transform 1 0 2162 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_282
timestamp 1571791925
transform 1 0 1334 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_283
timestamp 1571791925
transform 1 0 2346 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_284
timestamp 1571791925
transform 1 0 2530 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_285
timestamp 1571791925
transform 1 0 2162 0 1 3910
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_286
timestamp 1571791925
transform 1 0 1886 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_287
timestamp 1571791925
transform 1 0 2162 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_288
timestamp 1571791925
transform 1 0 2070 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_289
timestamp 1571791925
transform 1 0 2622 0 1 4182
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_290
timestamp 1571791925
transform 1 0 1426 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_291
timestamp 1571791925
transform 1 0 2990 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_292
timestamp 1571791925
transform 1 0 4830 0 1 4726
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_293
timestamp 1571791925
transform 1 0 4830 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_294
timestamp 1571791925
transform 1 0 3634 0 1 5202
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_295
timestamp 1571791925
transform 1 0 3818 0 1 2958
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_296
timestamp 1571791925
transform 1 0 4922 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_297
timestamp 1571791925
transform 1 0 3818 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_298
timestamp 1571791925
transform 1 0 4646 0 1 5134
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_299
timestamp 1571791925
transform 1 0 4646 0 1 4726
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_300
timestamp 1571791925
transform 1 0 4646 0 1 3570
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_301
timestamp 1571791925
transform 1 0 3450 0 1 3026
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_302
timestamp 1571791925
transform 1 0 4462 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_303
timestamp 1571791925
transform 1 0 4186 0 1 3094
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_304
timestamp 1571791925
transform 1 0 4094 0 1 3978
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_305
timestamp 1571791925
transform 1 0 4646 0 1 5270
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_306
timestamp 1571791925
transform 1 0 4646 0 1 4590
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_307
timestamp 1571791925
transform 1 0 3542 0 1 3502
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_308
timestamp 1571791925
transform 1 0 4830 0 1 3978
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_309
timestamp 1571791925
transform 1 0 4646 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_310
timestamp 1571791925
transform 1 0 3542 0 1 6970
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_311
timestamp 1571791925
transform 1 0 4186 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_312
timestamp 1571791925
transform 1 0 4646 0 1 6902
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_313
timestamp 1571791925
transform 1 0 4186 0 1 6902
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_314
timestamp 1571791925
transform 1 0 4278 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_315
timestamp 1571791925
transform 1 0 4278 0 1 6698
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_316
timestamp 1571791925
transform 1 0 3634 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_317
timestamp 1571791925
transform 1 0 4646 0 1 7922
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_318
timestamp 1571791925
transform 1 0 4830 0 1 6834
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_319
timestamp 1571791925
transform 1 0 4830 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_320
timestamp 1571791925
transform 1 0 4738 0 1 6630
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_321
timestamp 1571791925
transform 1 0 4738 0 1 7718
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_322
timestamp 1571791925
transform 1 0 4738 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_323
timestamp 1571791925
transform 1 0 1978 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_324
timestamp 1571791925
transform 1 0 2162 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_325
timestamp 1571791925
transform 1 0 2162 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_326
timestamp 1571791925
transform 1 0 2162 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_327
timestamp 1571791925
transform 1 0 2162 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_328
timestamp 1571791925
transform 1 0 1426 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_329
timestamp 1571791925
transform 1 0 1702 0 1 7922
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_330
timestamp 1571791925
transform 1 0 1426 0 1 6834
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_331
timestamp 1571791925
transform 1 0 2898 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_332
timestamp 1571791925
transform 1 0 1886 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_333
timestamp 1571791925
transform 1 0 2070 0 1 6698
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_334
timestamp 1571791925
transform 1 0 2070 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_335
timestamp 1571791925
transform 1 0 1426 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_336
timestamp 1571791925
transform 1 0 1978 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_337
timestamp 1571791925
transform 1 0 1886 0 1 9146
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_338
timestamp 1571791925
transform 1 0 1334 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_339
timestamp 1571791925
transform 1 0 1702 0 1 8330
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_340
timestamp 1571791925
transform 1 0 2162 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_341
timestamp 1571791925
transform 1 0 2162 0 1 9486
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_342
timestamp 1571791925
transform 1 0 1334 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_343
timestamp 1571791925
transform 1 0 2070 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_344
timestamp 1571791925
transform 1 0 2070 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_345
timestamp 1571791925
transform 1 0 3174 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_346
timestamp 1571791925
transform 1 0 2990 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_347
timestamp 1571791925
transform 1 0 2990 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_348
timestamp 1571791925
transform 1 0 3266 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_349
timestamp 1571791925
transform 1 0 3266 0 1 8058
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_350
timestamp 1571791925
transform 1 0 3266 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_351
timestamp 1571791925
transform 1 0 2990 0 1 8058
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_352
timestamp 1571791925
transform 1 0 1886 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_353
timestamp 1571791925
transform 1 0 2254 0 1 9010
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_354
timestamp 1571791925
transform 1 0 1978 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_355
timestamp 1571791925
transform 1 0 2254 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_356
timestamp 1571791925
transform 1 0 3910 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_357
timestamp 1571791925
transform 1 0 4738 0 1 9690
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_358
timestamp 1571791925
transform 1 0 4738 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_359
timestamp 1571791925
transform 1 0 4646 0 1 9010
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_360
timestamp 1571791925
transform 1 0 4186 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_361
timestamp 1571791925
transform 1 0 4186 0 1 9894
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_362
timestamp 1571791925
transform 1 0 4554 0 1 9350
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_363
timestamp 1571791925
transform 1 0 4646 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_364
timestamp 1571791925
transform 1 0 3910 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_365
timestamp 1571791925
transform 1 0 7958 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_366
timestamp 1571791925
transform 1 0 8326 0 1 6290
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_367
timestamp 1571791925
transform 1 0 8602 0 1 7446
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_368
timestamp 1571791925
transform 1 0 7682 0 1 7174
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_369
timestamp 1571791925
transform 1 0 7682 0 1 6698
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_370
timestamp 1571791925
transform 1 0 8050 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_371
timestamp 1571791925
transform 1 0 7774 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_372
timestamp 1571791925
transform 1 0 8602 0 1 6630
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_373
timestamp 1571791925
transform 1 0 8694 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_374
timestamp 1571791925
transform 1 0 8602 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_375
timestamp 1571791925
transform 1 0 8694 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_376
timestamp 1571791925
transform 1 0 7958 0 1 5746
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_377
timestamp 1571791925
transform 1 0 8234 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_378
timestamp 1571791925
transform 1 0 8510 0 1 5542
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_379
timestamp 1571791925
transform 1 0 8418 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_380
timestamp 1571791925
transform 1 0 8418 0 1 6834
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_381
timestamp 1571791925
transform 1 0 9338 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_382
timestamp 1571791925
transform 1 0 9338 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_383
timestamp 1571791925
transform 1 0 7498 0 1 6086
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_384
timestamp 1571791925
transform 1 0 8326 0 1 7310
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_385
timestamp 1571791925
transform 1 0 7958 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_386
timestamp 1571791925
transform 1 0 7038 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_387
timestamp 1571791925
transform 1 0 6486 0 1 7310
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_388
timestamp 1571791925
transform 1 0 5474 0 1 6698
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_389
timestamp 1571791925
transform 1 0 6486 0 1 6970
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_390
timestamp 1571791925
transform 1 0 5842 0 1 6086
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_391
timestamp 1571791925
transform 1 0 7038 0 1 6834
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_392
timestamp 1571791925
transform 1 0 5842 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_393
timestamp 1571791925
transform 1 0 6762 0 1 7446
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_394
timestamp 1571791925
transform 1 0 6486 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_395
timestamp 1571791925
transform 1 0 5658 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_396
timestamp 1571791925
transform 1 0 6854 0 1 5814
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_397
timestamp 1571791925
transform 1 0 6118 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_398
timestamp 1571791925
transform 1 0 6118 0 1 7718
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_399
timestamp 1571791925
transform 1 0 5566 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_400
timestamp 1571791925
transform 1 0 5566 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_401
timestamp 1571791925
transform 1 0 6946 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_402
timestamp 1571791925
transform 1 0 6302 0 1 6426
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_403
timestamp 1571791925
transform 1 0 5842 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_404
timestamp 1571791925
transform 1 0 5566 0 1 6222
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_405
timestamp 1571791925
transform 1 0 6394 0 1 5814
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_406
timestamp 1571791925
transform 1 0 7038 0 1 7514
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_407
timestamp 1571791925
transform 1 0 7406 0 1 7378
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_408
timestamp 1571791925
transform 1 0 5934 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_409
timestamp 1571791925
transform 1 0 5658 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_410
timestamp 1571791925
transform 1 0 5658 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_411
timestamp 1571791925
transform 1 0 5934 0 1 6358
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_412
timestamp 1571791925
transform 1 0 5750 0 1 7446
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_413
timestamp 1571791925
transform 1 0 5750 0 1 5678
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_414
timestamp 1571791925
transform 1 0 7406 0 1 6154
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_415
timestamp 1571791925
transform 1 0 5474 0 1 6154
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_416
timestamp 1571791925
transform 1 0 5934 0 1 7854
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_417
timestamp 1571791925
transform 1 0 6394 0 1 6766
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_418
timestamp 1571791925
transform 1 0 6762 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_419
timestamp 1571791925
transform 1 0 5474 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_420
timestamp 1571791925
transform 1 0 6486 0 1 9350
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_421
timestamp 1571791925
transform 1 0 5658 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_422
timestamp 1571791925
transform 1 0 5658 0 1 9146
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_423
timestamp 1571791925
transform 1 0 5474 0 1 10574
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_424
timestamp 1571791925
transform 1 0 5566 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_425
timestamp 1571791925
transform 1 0 6394 0 1 9146
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_426
timestamp 1571791925
transform 1 0 6394 0 1 9486
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_427
timestamp 1571791925
transform 1 0 6394 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_428
timestamp 1571791925
transform 1 0 6854 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_429
timestamp 1571791925
transform 1 0 6854 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_430
timestamp 1571791925
transform 1 0 7038 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_431
timestamp 1571791925
transform 1 0 6854 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_432
timestamp 1571791925
transform 1 0 5750 0 1 8806
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_433
timestamp 1571791925
transform 1 0 7130 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_434
timestamp 1571791925
transform 1 0 7038 0 1 9418
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_435
timestamp 1571791925
transform 1 0 6026 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_436
timestamp 1571791925
transform 1 0 6026 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_437
timestamp 1571791925
transform 1 0 7038 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_438
timestamp 1571791925
transform 1 0 5842 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_439
timestamp 1571791925
transform 1 0 5934 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_440
timestamp 1571791925
transform 1 0 9154 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_441
timestamp 1571791925
transform 1 0 9154 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_442
timestamp 1571791925
transform 1 0 8326 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_443
timestamp 1571791925
transform 1 0 8970 0 1 10234
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_444
timestamp 1571791925
transform 1 0 8326 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_445
timestamp 1571791925
transform 1 0 8326 0 1 8602
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_446
timestamp 1571791925
transform 1 0 9338 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_447
timestamp 1571791925
transform 1 0 7866 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_448
timestamp 1571791925
transform 1 0 9246 0 1 10098
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_449
timestamp 1571791925
transform 1 0 8326 0 1 10506
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_450
timestamp 1571791925
transform 1 0 8418 0 1 10030
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_451
timestamp 1571791925
transform 1 0 8510 0 1 8466
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_452
timestamp 1571791925
transform 1 0 8510 0 1 9486
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_453
timestamp 1571791925
transform 1 0 7866 0 1 9350
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_454
timestamp 1571791925
transform 1 0 7774 0 1 8534
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_455
timestamp 1571791925
transform 1 0 8970 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_456
timestamp 1571791925
transform 1 0 7774 0 1 9554
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_457
timestamp 1571791925
transform 1 0 9338 0 1 9622
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_458
timestamp 1571791925
transform 1 0 9246 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_459
timestamp 1571791925
transform 1 0 9246 0 1 8874
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_460
timestamp 1571791925
transform 1 0 8602 0 1 8942
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_461
timestamp 1571791925
transform 1 0 5750 0 1 7990
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_462
timestamp 1571791925
transform 1 0 5382 0 1 9962
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_463
timestamp 1571791925
transform 1 0 5382 0 1 4250
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_464
timestamp 1571791925
transform 1 0 5382 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_465
timestamp 1571791925
transform 1 0 6118 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_466
timestamp 1571791925
transform 1 0 5382 0 1 4114
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_467
timestamp 1571791925
transform 1 0 5382 0 1 7786
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_468
timestamp 1571791925
transform 1 0 5382 0 1 8398
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_469
timestamp 1571791925
transform 1 0 2898 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_470
timestamp 1571791925
transform 1 0 2346 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_471
timestamp 1571791925
transform 1 0 4738 0 1 5338
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_472
timestamp 1571791925
transform 1 0 8602 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_473
timestamp 1571791925
transform 1 0 9246 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_474
timestamp 1571791925
transform 1 0 9154 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_475
timestamp 1571791925
transform 1 0 7958 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_476
timestamp 1571791925
transform 1 0 7958 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_477
timestamp 1571791925
transform 1 0 9246 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_478
timestamp 1571791925
transform 1 0 7958 0 1 12886
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_479
timestamp 1571791925
transform 1 0 8970 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_480
timestamp 1571791925
transform 1 0 9062 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_481
timestamp 1571791925
transform 1 0 9338 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_482
timestamp 1571791925
transform 1 0 8418 0 1 11322
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_483
timestamp 1571791925
transform 1 0 9154 0 1 10982
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_484
timestamp 1571791925
transform 1 0 8326 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_485
timestamp 1571791925
transform 1 0 8602 0 1 12886
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_486
timestamp 1571791925
transform 1 0 7866 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_487
timestamp 1571791925
transform 1 0 7866 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_488
timestamp 1571791925
transform 1 0 8418 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_489
timestamp 1571791925
transform 1 0 9246 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_490
timestamp 1571791925
transform 1 0 6854 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_491
timestamp 1571791925
transform 1 0 5934 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_492
timestamp 1571791925
transform 1 0 5842 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_493
timestamp 1571791925
transform 1 0 5750 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_494
timestamp 1571791925
transform 1 0 6946 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_495
timestamp 1571791925
transform 1 0 5750 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_496
timestamp 1571791925
transform 1 0 5474 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_497
timestamp 1571791925
transform 1 0 6762 0 1 12274
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_498
timestamp 1571791925
transform 1 0 6946 0 1 12614
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_499
timestamp 1571791925
transform 1 0 6762 0 1 11322
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_500
timestamp 1571791925
transform 1 0 6394 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_501
timestamp 1571791925
transform 1 0 6854 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_502
timestamp 1571791925
transform 1 0 7130 0 1 10710
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_503
timestamp 1571791925
transform 1 0 5566 0 1 10982
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_504
timestamp 1571791925
transform 1 0 6118 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_505
timestamp 1571791925
transform 1 0 5934 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_506
timestamp 1571791925
transform 1 0 5842 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_507
timestamp 1571791925
transform 1 0 7038 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_508
timestamp 1571791925
transform 1 0 6670 0 1 12954
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_509
timestamp 1571791925
transform 1 0 6394 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_510
timestamp 1571791925
transform 1 0 7314 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_511
timestamp 1571791925
transform 1 0 5750 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_512
timestamp 1571791925
transform 1 0 6302 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_513
timestamp 1571791925
transform 1 0 6302 0 1 14042
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_514
timestamp 1571791925
transform 1 0 5842 0 1 13974
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_515
timestamp 1571791925
transform 1 0 7038 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_516
timestamp 1571791925
transform 1 0 5842 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_517
timestamp 1571791925
transform 1 0 6118 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_518
timestamp 1571791925
transform 1 0 6118 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_519
timestamp 1571791925
transform 1 0 5750 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_520
timestamp 1571791925
transform 1 0 5750 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_521
timestamp 1571791925
transform 1 0 7314 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_522
timestamp 1571791925
transform 1 0 7406 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_523
timestamp 1571791925
transform 1 0 6946 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_524
timestamp 1571791925
transform 1 0 6946 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_525
timestamp 1571791925
transform 1 0 7222 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_526
timestamp 1571791925
transform 1 0 7038 0 1 14518
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_527
timestamp 1571791925
transform 1 0 6670 0 1 15674
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_528
timestamp 1571791925
transform 1 0 7406 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_529
timestamp 1571791925
transform 1 0 6670 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_530
timestamp 1571791925
transform 1 0 7222 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_531
timestamp 1571791925
transform 1 0 5474 0 1 13362
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_532
timestamp 1571791925
transform 1 0 6670 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_533
timestamp 1571791925
transform 1 0 6670 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_534
timestamp 1571791925
transform 1 0 9246 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_535
timestamp 1571791925
transform 1 0 7590 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_536
timestamp 1571791925
transform 1 0 7590 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_537
timestamp 1571791925
transform 1 0 7590 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_538
timestamp 1571791925
transform 1 0 7590 0 1 14790
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_539
timestamp 1571791925
transform 1 0 9154 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_540
timestamp 1571791925
transform 1 0 9246 0 1 13974
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_541
timestamp 1571791925
transform 1 0 9246 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_542
timestamp 1571791925
transform 1 0 8786 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_543
timestamp 1571791925
transform 1 0 8786 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_544
timestamp 1571791925
transform 1 0 8510 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_545
timestamp 1571791925
transform 1 0 8510 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_546
timestamp 1571791925
transform 1 0 7958 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_547
timestamp 1571791925
transform 1 0 7682 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_548
timestamp 1571791925
transform 1 0 8326 0 1 13362
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_549
timestamp 1571791925
transform 1 0 7682 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_550
timestamp 1571791925
transform 1 0 9338 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_551
timestamp 1571791925
transform 1 0 9338 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_552
timestamp 1571791925
transform 1 0 9154 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_553
timestamp 1571791925
transform 1 0 6946 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_554
timestamp 1571791925
transform 1 0 4646 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_555
timestamp 1571791925
transform 1 0 3818 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_556
timestamp 1571791925
transform 1 0 3818 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_557
timestamp 1571791925
transform 1 0 5290 0 1 11798
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_558
timestamp 1571791925
transform 1 0 4094 0 1 11594
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_559
timestamp 1571791925
transform 1 0 4738 0 1 11322
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_560
timestamp 1571791925
transform 1 0 4738 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_561
timestamp 1571791925
transform 1 0 4002 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_562
timestamp 1571791925
transform 1 0 4002 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_563
timestamp 1571791925
transform 1 0 3542 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_564
timestamp 1571791925
transform 1 0 3542 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_565
timestamp 1571791925
transform 1 0 4646 0 1 12954
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_566
timestamp 1571791925
transform 1 0 4830 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_567
timestamp 1571791925
transform 1 0 3450 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_568
timestamp 1571791925
transform 1 0 4830 0 1 10710
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_569
timestamp 1571791925
transform 1 0 4646 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_570
timestamp 1571791925
transform 1 0 5198 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_571
timestamp 1571791925
transform 1 0 5198 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_572
timestamp 1571791925
transform 1 0 4830 0 1 12614
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_573
timestamp 1571791925
transform 1 0 4094 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_574
timestamp 1571791925
transform 1 0 4738 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_575
timestamp 1571791925
transform 1 0 1426 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_576
timestamp 1571791925
transform 1 0 3174 0 1 11322
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_577
timestamp 1571791925
transform 1 0 3174 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_578
timestamp 1571791925
transform 1 0 1518 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_579
timestamp 1571791925
transform 1 0 2254 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_580
timestamp 1571791925
transform 1 0 1518 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_581
timestamp 1571791925
transform 1 0 1426 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_582
timestamp 1571791925
transform 1 0 1794 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_583
timestamp 1571791925
transform 1 0 1794 0 1 10710
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_584
timestamp 1571791925
transform 1 0 2254 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_585
timestamp 1571791925
transform 1 0 2070 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_586
timestamp 1571791925
transform 1 0 2070 0 1 12070
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_587
timestamp 1571791925
transform 1 0 2806 0 1 12274
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_588
timestamp 1571791925
transform 1 0 1978 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_589
timestamp 1571791925
transform 1 0 1978 0 1 10710
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_590
timestamp 1571791925
transform 1 0 2162 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_591
timestamp 1571791925
transform 1 0 2806 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_592
timestamp 1571791925
transform 1 0 2162 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_593
timestamp 1571791925
transform 1 0 2806 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_594
timestamp 1571791925
transform 1 0 2806 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_595
timestamp 1571791925
transform 1 0 2346 0 1 14790
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_596
timestamp 1571791925
transform 1 0 2346 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_597
timestamp 1571791925
transform 1 0 2806 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_598
timestamp 1571791925
transform 1 0 1978 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_599
timestamp 1571791925
transform 1 0 1978 0 1 13974
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_600
timestamp 1571791925
transform 1 0 2070 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_601
timestamp 1571791925
transform 1 0 1978 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_602
timestamp 1571791925
transform 1 0 2070 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_603
timestamp 1571791925
transform 1 0 1426 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_604
timestamp 1571791925
transform 1 0 1334 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_605
timestamp 1571791925
transform 1 0 1334 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_606
timestamp 1571791925
transform 1 0 3174 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_607
timestamp 1571791925
transform 1 0 3174 0 1 13498
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_608
timestamp 1571791925
transform 1 0 2806 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_609
timestamp 1571791925
transform 1 0 2254 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_610
timestamp 1571791925
transform 1 0 2898 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_611
timestamp 1571791925
transform 1 0 2898 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_612
timestamp 1571791925
transform 1 0 1702 0 1 13362
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_613
timestamp 1571791925
transform 1 0 1702 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_614
timestamp 1571791925
transform 1 0 1794 0 1 15538
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_615
timestamp 1571791925
transform 1 0 2070 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_616
timestamp 1571791925
transform 1 0 4094 0 1 15538
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_617
timestamp 1571791925
transform 1 0 4646 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_618
timestamp 1571791925
transform 1 0 4646 0 1 13362
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_619
timestamp 1571791925
transform 1 0 3542 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_620
timestamp 1571791925
transform 1 0 4646 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_621
timestamp 1571791925
transform 1 0 4738 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_622
timestamp 1571791925
transform 1 0 5014 0 1 15538
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_623
timestamp 1571791925
transform 1 0 4186 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_624
timestamp 1571791925
transform 1 0 3542 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_625
timestamp 1571791925
transform 1 0 4002 0 1 15674
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_626
timestamp 1571791925
transform 1 0 4646 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_627
timestamp 1571791925
transform 1 0 3358 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_628
timestamp 1571791925
transform 1 0 3358 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_629
timestamp 1571791925
transform 1 0 3358 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_630
timestamp 1571791925
transform 1 0 3358 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_631
timestamp 1571791925
transform 1 0 4002 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_632
timestamp 1571791925
transform 1 0 4094 0 1 16014
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_633
timestamp 1571791925
transform 1 0 4646 0 1 16490
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_634
timestamp 1571791925
transform 1 0 4186 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_635
timestamp 1571791925
transform 1 0 4186 0 1 16422
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_636
timestamp 1571791925
transform 1 0 4646 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_637
timestamp 1571791925
transform 1 0 4830 0 1 18394
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_638
timestamp 1571791925
transform 1 0 4830 0 1 17646
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_639
timestamp 1571791925
transform 1 0 3818 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_640
timestamp 1571791925
transform 1 0 3634 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_641
timestamp 1571791925
transform 1 0 3634 0 1 18326
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_642
timestamp 1571791925
transform 1 0 3818 0 1 16694
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_643
timestamp 1571791925
transform 1 0 4646 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_644
timestamp 1571791925
transform 1 0 3634 0 1 17714
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_645
timestamp 1571791925
transform 1 0 4002 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_646
timestamp 1571791925
transform 1 0 5014 0 1 16014
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_647
timestamp 1571791925
transform 1 0 3266 0 1 16422
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_648
timestamp 1571791925
transform 1 0 1702 0 1 16490
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_649
timestamp 1571791925
transform 1 0 1518 0 1 18258
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_650
timestamp 1571791925
transform 1 0 2346 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_651
timestamp 1571791925
transform 1 0 1610 0 1 18054
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_652
timestamp 1571791925
transform 1 0 3174 0 1 18054
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_653
timestamp 1571791925
transform 1 0 1518 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_654
timestamp 1571791925
transform 1 0 2990 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_655
timestamp 1571791925
transform 1 0 2990 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_656
timestamp 1571791925
transform 1 0 2990 0 1 17170
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_657
timestamp 1571791925
transform 1 0 1978 0 1 18258
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_658
timestamp 1571791925
transform 1 0 2990 0 1 18190
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_659
timestamp 1571791925
transform 1 0 1610 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_660
timestamp 1571791925
transform 1 0 2162 0 1 16490
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_661
timestamp 1571791925
transform 1 0 2254 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_662
timestamp 1571791925
transform 1 0 2806 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_663
timestamp 1571791925
transform 1 0 1794 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_664
timestamp 1571791925
transform 1 0 1794 0 1 17714
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_665
timestamp 1571791925
transform 1 0 3174 0 1 17850
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_666
timestamp 1571791925
transform 1 0 3266 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_667
timestamp 1571791925
transform 1 0 2898 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_668
timestamp 1571791925
transform 1 0 2162 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_669
timestamp 1571791925
transform 1 0 2806 0 1 17850
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_670
timestamp 1571791925
transform 1 0 1702 0 1 16150
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_671
timestamp 1571791925
transform 1 0 1978 0 1 18666
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_672
timestamp 1571791925
transform 1 0 2254 0 1 18734
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_673
timestamp 1571791925
transform 1 0 4738 0 1 18666
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_674
timestamp 1571791925
transform 1 0 4646 0 1 18598
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_675
timestamp 1571791925
transform 1 0 3818 0 1 18666
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_676
timestamp 1571791925
transform 1 0 4830 0 1 18734
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_677
timestamp 1571791925
transform 1 0 3358 0 1 18190
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_678
timestamp 1571791925
transform 1 0 3358 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_679
timestamp 1571791925
transform 1 0 8786 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_680
timestamp 1571791925
transform 1 0 8878 0 1 16014
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_681
timestamp 1571791925
transform 1 0 6210 0 1 18258
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_682
timestamp 1571791925
transform 1 0 6210 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_683
timestamp 1571791925
transform 1 0 5658 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_684
timestamp 1571791925
transform 1 0 5658 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_685
timestamp 1571791925
transform 1 0 5750 0 1 18258
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_686
timestamp 1571791925
transform 1 0 9338 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_687
timestamp 1571791925
transform 1 0 9338 0 1 16966
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_688
timestamp 1571791925
transform 1 0 9246 0 1 17170
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_689
timestamp 1571791925
transform 1 0 9246 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_690
timestamp 1571791925
transform 1 0 5474 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_691
timestamp 1571791925
transform 1 0 5474 0 1 18394
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_692
timestamp 1571791925
transform 1 0 7590 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_693
timestamp 1571791925
transform 1 0 7498 0 1 18734
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_694
timestamp 1571791925
transform 1 0 7498 0 1 18258
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_695
timestamp 1571791925
transform 1 0 7130 0 1 16966
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_696
timestamp 1571791925
transform 1 0 9338 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_697
timestamp 1571791925
transform 1 0 9338 0 1 17170
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_698
timestamp 1571791925
transform 1 0 5566 0 1 18326
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_699
timestamp 1571791925
transform 1 0 5566 0 1 16694
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_700
timestamp 1571791925
transform 1 0 7406 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_701
timestamp 1571791925
transform 1 0 7130 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_702
timestamp 1571791925
transform 1 0 9430 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_703
timestamp 1571791925
transform 1 0 7774 0 1 17646
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_704
timestamp 1571791925
transform 1 0 7774 0 1 18054
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_705
timestamp 1571791925
transform 1 0 9430 0 1 16490
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_706
timestamp 1571791925
transform 1 0 9430 0 1 18190
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_707
timestamp 1571791925
transform 1 0 9430 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_708
timestamp 1571791925
transform 1 0 6670 0 1 17714
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_709
timestamp 1571791925
transform 1 0 8786 0 1 17782
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_710
timestamp 1571791925
transform 1 0 6670 0 1 17102
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_711
timestamp 1571791925
transform 1 0 8786 0 1 18190
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_712
timestamp 1571791925
transform 1 0 5658 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_713
timestamp 1571791925
transform 1 0 5658 0 1 18122
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_714
timestamp 1571791925
transform 1 0 8234 0 1 18598
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_715
timestamp 1571791925
transform 1 0 6486 0 1 17646
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_716
timestamp 1571791925
transform 1 0 6486 0 1 18054
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_717
timestamp 1571791925
transform 1 0 7774 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_718
timestamp 1571791925
transform 1 0 5750 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_719
timestamp 1571791925
transform 1 0 7774 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_720
timestamp 1571791925
transform 1 0 7038 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_721
timestamp 1571791925
transform 1 0 7038 0 1 17102
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_722
timestamp 1571791925
transform 1 0 6118 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_723
timestamp 1571791925
transform 1 0 7682 0 1 17102
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_724
timestamp 1571791925
transform 1 0 8510 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_725
timestamp 1571791925
transform 1 0 8510 0 1 17646
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_726
timestamp 1571791925
transform 1 0 6026 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_727
timestamp 1571791925
transform 1 0 8234 0 1 18326
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_728
timestamp 1571791925
transform 1 0 6762 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_729
timestamp 1571791925
transform 1 0 6118 0 1 17170
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_730
timestamp 1571791925
transform 1 0 6762 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_731
timestamp 1571791925
transform 1 0 5382 0 1 15674
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_732
timestamp 1571791925
transform 1 0 5382 0 1 15878
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_733
timestamp 1571791925
transform 1 0 5382 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_734
timestamp 1571791925
transform 1 0 5382 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_735
timestamp 1571791925
transform 1 0 5382 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_736
timestamp 1571791925
transform 1 0 17342 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_737
timestamp 1571791925
transform 1 0 17342 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_738
timestamp 1571791925
transform 1 0 16606 0 1 12614
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_739
timestamp 1571791925
transform 1 0 16606 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_740
timestamp 1571791925
transform 1 0 17066 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_741
timestamp 1571791925
transform 1 0 17342 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_742
timestamp 1571791925
transform 1 0 16882 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_743
timestamp 1571791925
transform 1 0 17066 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_744
timestamp 1571791925
transform 1 0 16882 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_745
timestamp 1571791925
transform 1 0 17434 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_746
timestamp 1571791925
transform 1 0 17526 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_747
timestamp 1571791925
transform 1 0 15778 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_748
timestamp 1571791925
transform 1 0 14490 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_749
timestamp 1571791925
transform 1 0 14490 0 1 12274
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_750
timestamp 1571791925
transform 1 0 13846 0 1 12682
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_751
timestamp 1571791925
transform 1 0 15410 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_752
timestamp 1571791925
transform 1 0 14490 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_753
timestamp 1571791925
transform 1 0 14490 0 1 11526
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_754
timestamp 1571791925
transform 1 0 14122 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_755
timestamp 1571791925
transform 1 0 14766 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_756
timestamp 1571791925
transform 1 0 14766 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_757
timestamp 1571791925
transform 1 0 14122 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_758
timestamp 1571791925
transform 1 0 15410 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_759
timestamp 1571791925
transform 1 0 14214 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_760
timestamp 1571791925
transform 1 0 14214 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_761
timestamp 1571791925
transform 1 0 14214 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_762
timestamp 1571791925
transform 1 0 14858 0 1 11186
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_763
timestamp 1571791925
transform 1 0 14858 0 1 11594
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_764
timestamp 1571791925
transform 1 0 13662 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_765
timestamp 1571791925
transform 1 0 15410 0 1 12274
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_766
timestamp 1571791925
transform 1 0 13662 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_767
timestamp 1571791925
transform 1 0 15318 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_768
timestamp 1571791925
transform 1 0 14950 0 1 12274
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_769
timestamp 1571791925
transform 1 0 14950 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_770
timestamp 1571791925
transform 1 0 15502 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_771
timestamp 1571791925
transform 1 0 15502 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_772
timestamp 1571791925
transform 1 0 13846 0 1 13362
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_773
timestamp 1571791925
transform 1 0 15226 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_774
timestamp 1571791925
transform 1 0 15226 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_775
timestamp 1571791925
transform 1 0 14674 0 1 14790
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_776
timestamp 1571791925
transform 1 0 14766 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_777
timestamp 1571791925
transform 1 0 14674 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_778
timestamp 1571791925
transform 1 0 15410 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_779
timestamp 1571791925
transform 1 0 15318 0 1 13430
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_780
timestamp 1571791925
transform 1 0 15502 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_781
timestamp 1571791925
transform 1 0 15502 0 1 14586
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_782
timestamp 1571791925
transform 1 0 15410 0 1 13974
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_783
timestamp 1571791925
transform 1 0 14214 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_784
timestamp 1571791925
transform 1 0 14214 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_785
timestamp 1571791925
transform 1 0 15594 0 1 15130
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_786
timestamp 1571791925
transform 1 0 15594 0 1 13498
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_787
timestamp 1571791925
transform 1 0 14398 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_788
timestamp 1571791925
transform 1 0 14398 0 1 14858
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_789
timestamp 1571791925
transform 1 0 14306 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_790
timestamp 1571791925
transform 1 0 15778 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_791
timestamp 1571791925
transform 1 0 15870 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_792
timestamp 1571791925
transform 1 0 15870 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_793
timestamp 1571791925
transform 1 0 15686 0 1 14790
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_794
timestamp 1571791925
transform 1 0 15686 0 1 12886
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_795
timestamp 1571791925
transform 1 0 15686 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_796
timestamp 1571791925
transform 1 0 15686 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_797
timestamp 1571791925
transform 1 0 15686 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_798
timestamp 1571791925
transform 1 0 15686 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_799
timestamp 1571791925
transform 1 0 15870 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_800
timestamp 1571791925
transform 1 0 12374 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_801
timestamp 1571791925
transform 1 0 12374 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_802
timestamp 1571791925
transform 1 0 12190 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_803
timestamp 1571791925
transform 1 0 13386 0 1 12750
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_804
timestamp 1571791925
transform 1 0 13386 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_805
timestamp 1571791925
transform 1 0 12558 0 1 11730
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_806
timestamp 1571791925
transform 1 0 12558 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_807
timestamp 1571791925
transform 1 0 13018 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_808
timestamp 1571791925
transform 1 0 12926 0 1 10710
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_809
timestamp 1571791925
transform 1 0 12926 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_810
timestamp 1571791925
transform 1 0 12098 0 1 11866
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_811
timestamp 1571791925
transform 1 0 12098 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_812
timestamp 1571791925
transform 1 0 12834 0 1 12070
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_813
timestamp 1571791925
transform 1 0 12006 0 1 10982
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_814
timestamp 1571791925
transform 1 0 12834 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_815
timestamp 1571791925
transform 1 0 11638 0 1 12138
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_816
timestamp 1571791925
transform 1 0 12466 0 1 13158
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_817
timestamp 1571791925
transform 1 0 12466 0 1 12342
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_818
timestamp 1571791925
transform 1 0 11822 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_819
timestamp 1571791925
transform 1 0 11822 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_820
timestamp 1571791925
transform 1 0 13386 0 1 11662
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_821
timestamp 1571791925
transform 1 0 13386 0 1 11118
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_822
timestamp 1571791925
transform 1 0 9706 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_823
timestamp 1571791925
transform 1 0 9798 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_824
timestamp 1571791925
transform 1 0 10074 0 1 12206
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_825
timestamp 1571791925
transform 1 0 10074 0 1 12682
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_826
timestamp 1571791925
transform 1 0 10626 0 1 12410
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_827
timestamp 1571791925
transform 1 0 10718 0 1 10778
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_828
timestamp 1571791925
transform 1 0 10718 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_829
timestamp 1571791925
transform 1 0 9982 0 1 11050
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_830
timestamp 1571791925
transform 1 0 10810 0 1 10642
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_831
timestamp 1571791925
transform 1 0 11362 0 1 12070
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_832
timestamp 1571791925
transform 1 0 9706 0 1 12818
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_833
timestamp 1571791925
transform 1 0 11454 0 1 14246
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_834
timestamp 1571791925
transform 1 0 10074 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_835
timestamp 1571791925
transform 1 0 10074 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_836
timestamp 1571791925
transform 1 0 11454 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_837
timestamp 1571791925
transform 1 0 11362 0 1 14858
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_838
timestamp 1571791925
transform 1 0 11086 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_839
timestamp 1571791925
transform 1 0 11086 0 1 14858
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_840
timestamp 1571791925
transform 1 0 10258 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_841
timestamp 1571791925
transform 1 0 10258 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_842
timestamp 1571791925
transform 1 0 11270 0 1 14790
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_843
timestamp 1571791925
transform 1 0 11270 0 1 14314
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_844
timestamp 1571791925
transform 1 0 10810 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_845
timestamp 1571791925
transform 1 0 10810 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_846
timestamp 1571791925
transform 1 0 11178 0 1 13294
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_847
timestamp 1571791925
transform 1 0 11178 0 1 13498
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_848
timestamp 1571791925
transform 1 0 12834 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_849
timestamp 1571791925
transform 1 0 12834 0 1 14586
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_850
timestamp 1571791925
transform 1 0 12006 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_851
timestamp 1571791925
transform 1 0 12006 0 1 14586
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_852
timestamp 1571791925
transform 1 0 12190 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_853
timestamp 1571791925
transform 1 0 12190 0 1 15470
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_854
timestamp 1571791925
transform 1 0 11822 0 1 15606
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_855
timestamp 1571791925
transform 1 0 12742 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_856
timestamp 1571791925
transform 1 0 12742 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_857
timestamp 1571791925
transform 1 0 11638 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_858
timestamp 1571791925
transform 1 0 11822 0 1 14994
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_859
timestamp 1571791925
transform 1 0 11822 0 1 13906
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_860
timestamp 1571791925
transform 1 0 12834 0 1 13498
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_861
timestamp 1571791925
transform 1 0 13018 0 1 13498
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_862
timestamp 1571791925
transform 1 0 11822 0 1 15402
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_863
timestamp 1571791925
transform 1 0 13018 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_864
timestamp 1571791925
transform 1 0 13018 0 1 15606
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_865
timestamp 1571791925
transform 1 0 13110 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_866
timestamp 1571791925
transform 1 0 12466 0 1 14382
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_867
timestamp 1571791925
transform 1 0 12466 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_868
timestamp 1571791925
transform 1 0 13202 0 1 15062
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_869
timestamp 1571791925
transform 1 0 13202 0 1 15334
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_870
timestamp 1571791925
transform 1 0 12558 0 1 14450
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_871
timestamp 1571791925
transform 1 0 12558 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_872
timestamp 1571791925
transform 1 0 12926 0 1 14926
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_873
timestamp 1571791925
transform 1 0 12926 0 1 14518
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_874
timestamp 1571791925
transform 1 0 13294 0 1 13702
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_875
timestamp 1571791925
transform 1 0 11638 0 1 13838
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_876
timestamp 1571791925
transform 1 0 12190 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_877
timestamp 1571791925
transform 1 0 9798 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_878
timestamp 1571791925
transform 1 0 11270 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_879
timestamp 1571791925
transform 1 0 11546 0 1 12886
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_880
timestamp 1571791925
transform 1 0 13294 0 1 13226
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_881
timestamp 1571791925
transform 1 0 10534 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_882
timestamp 1571791925
transform 1 0 10534 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_883
timestamp 1571791925
transform 1 0 11362 0 1 17646
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_884
timestamp 1571791925
transform 1 0 11362 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_885
timestamp 1571791925
transform 1 0 12006 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_886
timestamp 1571791925
transform 1 0 12006 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_887
timestamp 1571791925
transform 1 0 10626 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_888
timestamp 1571791925
transform 1 0 10810 0 1 17170
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_889
timestamp 1571791925
transform 1 0 10074 0 1 18734
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_890
timestamp 1571791925
transform 1 0 10810 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_891
timestamp 1571791925
transform 1 0 10810 0 1 16558
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_892
timestamp 1571791925
transform 1 0 10074 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_893
timestamp 1571791925
transform 1 0 11822 0 1 16966
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_894
timestamp 1571791925
transform 1 0 13110 0 1 16966
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_895
timestamp 1571791925
transform 1 0 10718 0 1 16762
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_896
timestamp 1571791925
transform 1 0 10718 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_897
timestamp 1571791925
transform 1 0 11822 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_898
timestamp 1571791925
transform 1 0 11822 0 1 17510
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_899
timestamp 1571791925
transform 1 0 11178 0 1 18054
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_900
timestamp 1571791925
transform 1 0 11178 0 1 17714
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_901
timestamp 1571791925
transform 1 0 11362 0 1 17102
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_902
timestamp 1571791925
transform 1 0 11362 0 1 16694
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_903
timestamp 1571791925
transform 1 0 9706 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_904
timestamp 1571791925
transform 1 0 9706 0 1 18190
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_905
timestamp 1571791925
transform 1 0 11546 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_906
timestamp 1571791925
transform 1 0 11362 0 1 16082
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_907
timestamp 1571791925
transform 1 0 10166 0 1 16218
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_908
timestamp 1571791925
transform 1 0 10166 0 1 16490
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_909
timestamp 1571791925
transform 1 0 10442 0 1 18326
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_910
timestamp 1571791925
transform 1 0 10442 0 1 18598
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_911
timestamp 1571791925
transform 1 0 12558 0 1 16762
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_912
timestamp 1571791925
transform 1 0 12558 0 1 17238
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_913
timestamp 1571791925
transform 1 0 14306 0 1 16626
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_914
timestamp 1571791925
transform 1 0 12926 0 1 15878
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_915
timestamp 1571791925
transform 1 0 9522 0 1 5610
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_916
timestamp 1571791925
transform 1 0 9522 0 1 4794
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_917
timestamp 1571791925
transform 1 0 9522 0 1 17578
box -32 -32 32 32
use VIA_M1M2_PR  VIA_M1M2_PR_918
timestamp 1571791925
transform 1 0 9522 0 1 17306
box -32 -32 32 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_0
timestamp 1571791925
transform 1 0 16606 0 1 8942
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_1
timestamp 1571791925
transform 1 0 4738 0 1 5678
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_2
timestamp 1571791925
transform 1 0 4738 0 1 10030
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_3
timestamp 1571791925
transform 1 0 8326 0 1 11730
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_4
timestamp 1571791925
transform 1 0 4738 0 1 17646
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_5
timestamp 1571791925
transform 1 0 6026 0 1 17170
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_6
timestamp 1571791925
transform 1 0 16606 0 1 11118
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_7
timestamp 1571791925
transform 1 0 12006 0 1 10642
box -26 -32 26 32
use VIA_M1M2_PR_MR  VIA_M1M2_PR_MR_8
timestamp 1571791925
transform 1 0 10626 0 1 12818
box -26 -32 26 32
use VIA_M2M3_PR  VIA_M2M3_PR_0
timestamp 1571791925
transform 1 0 12466 0 1 748
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_1
timestamp 1571791925
transform 1 0 12834 0 1 68
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_2
timestamp 1571791925
transform 1 0 10350 0 1 6868
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_3
timestamp 1571791925
transform 1 0 10350 0 1 6188
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_4
timestamp 1571791925
transform 1 0 17158 0 1 9588
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_5
timestamp 1571791925
transform 1 0 15870 0 1 10540
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_6
timestamp 1571791925
transform 1 0 8970 0 1 1428
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_7
timestamp 1571791925
transform 1 0 6394 0 1 2380
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_8
timestamp 1571791925
transform 1 0 5934 0 1 5100
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_9
timestamp 1571791925
transform 1 0 7682 0 1 5236
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_10
timestamp 1571791925
transform 1 0 8326 0 1 5236
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_11
timestamp 1571791925
transform 1 0 1334 0 1 4148
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_12
timestamp 1571791925
transform 1 0 2162 0 1 2788
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_13
timestamp 1571791925
transform 1 0 1702 0 1 2788
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_14
timestamp 1571791925
transform 1 0 4922 0 1 3468
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_15
timestamp 1571791925
transform 1 0 1334 0 1 8908
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_16
timestamp 1571791925
transform 1 0 4646 0 1 9588
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_17
timestamp 1571791925
transform 1 0 4738 0 1 7956
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_18
timestamp 1571791925
transform 1 0 7774 0 1 7820
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_19
timestamp 1571791925
transform 1 0 5474 0 1 9588
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_20
timestamp 1571791925
transform 1 0 8970 0 1 10132
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_21
timestamp 1571791925
transform 1 0 9246 0 1 12852
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_22
timestamp 1571791925
transform 1 0 7314 0 1 13396
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_23
timestamp 1571791925
transform 1 0 1518 0 1 11628
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_24
timestamp 1571791925
transform 1 0 1334 0 1 15028
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_25
timestamp 1571791925
transform 1 0 2898 0 1 15708
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_26
timestamp 1571791925
transform 1 0 4186 0 1 14348
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_27
timestamp 1571791925
transform 1 0 4554 0 1 16388
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_28
timestamp 1571791925
transform 1 0 2254 0 1 19108
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_29
timestamp 1571791925
transform 1 0 2806 0 1 20468
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_30
timestamp 1571791925
transform 1 0 1518 0 1 19788
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_31
timestamp 1571791925
transform 1 0 3450 0 1 21148
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_32
timestamp 1571791925
transform 1 0 9246 0 1 17068
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_33
timestamp 1571791925
transform 1 0 17526 0 1 10948
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_34
timestamp 1571791925
transform 1 0 17066 0 1 11628
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_35
timestamp 1571791925
transform 1 0 17618 0 1 11628
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_36
timestamp 1571791925
transform 1 0 11822 0 1 10676
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_37
timestamp 1571791925
transform 1 0 11362 0 1 12308
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_38
timestamp 1571791925
transform 1 0 10626 0 1 17748
box -33 -37 33 37
use VIA_M2M3_PR  VIA_M2M3_PR_39
timestamp 1571791925
transform 1 0 11638 0 1 18292
box -33 -37 33 37
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_0
timestamp 1571791925
transform 1 0 16368 0 1 3808
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_1
timestamp 1571791925
transform 1 0 17108 0 1 2176
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_2
timestamp 1571791925
transform 1 0 17108 0 1 4352
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_3
timestamp 1571791925
transform 1 0 16368 0 1 2720
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_4
timestamp 1571791925
transform 1 0 17108 0 1 3264
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_5
timestamp 1571791925
transform 1 0 16368 0 1 4896
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_6
timestamp 1571791925
transform 1 0 11108 0 1 2176
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_7
timestamp 1571791925
transform 1 0 10368 0 1 3808
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_8
timestamp 1571791925
transform 1 0 11108 0 1 3264
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_9
timestamp 1571791925
transform 1 0 11108 0 1 4352
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_10
timestamp 1571791925
transform 1 0 10368 0 1 4896
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_11
timestamp 1571791925
transform 1 0 10368 0 1 2720
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_12
timestamp 1571791925
transform 1 0 11108 0 1 7616
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_13
timestamp 1571791925
transform 1 0 10368 0 1 5984
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_14
timestamp 1571791925
transform 1 0 11108 0 1 5440
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_15
timestamp 1571791925
transform 1 0 10368 0 1 7072
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_16
timestamp 1571791925
transform 1 0 11108 0 1 6528
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_17
timestamp 1571791925
transform 1 0 11108 0 1 9792
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_18
timestamp 1571791925
transform 1 0 10368 0 1 10336
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_19
timestamp 1571791925
transform 1 0 10368 0 1 9248
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_20
timestamp 1571791925
transform 1 0 10368 0 1 8160
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_21
timestamp 1571791925
transform 1 0 11108 0 1 8704
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_22
timestamp 1571791925
transform 1 0 17108 0 1 5440
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_23
timestamp 1571791925
transform 1 0 16368 0 1 5984
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_24
timestamp 1571791925
transform 1 0 17108 0 1 7616
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_25
timestamp 1571791925
transform 1 0 17108 0 1 6528
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_26
timestamp 1571791925
transform 1 0 16368 0 1 7072
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_27
timestamp 1571791925
transform 1 0 16368 0 1 10336
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_28
timestamp 1571791925
transform 1 0 16368 0 1 8160
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_29
timestamp 1571791925
transform 1 0 16368 0 1 9248
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_30
timestamp 1571791925
transform 1 0 17108 0 1 9792
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_31
timestamp 1571791925
transform 1 0 17108 0 1 8704
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_32
timestamp 1571791925
transform 1 0 5108 0 1 2176
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_33
timestamp 1571791925
transform 1 0 4368 0 1 3808
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_34
timestamp 1571791925
transform 1 0 4368 0 1 4896
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_35
timestamp 1571791925
transform 1 0 5108 0 1 4352
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_36
timestamp 1571791925
transform 1 0 5108 0 1 3264
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_37
timestamp 1571791925
transform 1 0 4368 0 1 2720
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_38
timestamp 1571791925
transform 1 0 5108 0 1 6528
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_39
timestamp 1571791925
transform 1 0 5108 0 1 5440
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_40
timestamp 1571791925
transform 1 0 4368 0 1 7072
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_41
timestamp 1571791925
transform 1 0 5108 0 1 7616
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_42
timestamp 1571791925
transform 1 0 4368 0 1 5984
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_43
timestamp 1571791925
transform 1 0 5108 0 1 9792
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_44
timestamp 1571791925
transform 1 0 5108 0 1 8704
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_45
timestamp 1571791925
transform 1 0 4368 0 1 9248
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_46
timestamp 1571791925
transform 1 0 4368 0 1 10336
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_47
timestamp 1571791925
transform 1 0 4368 0 1 8160
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_48
timestamp 1571791925
transform 1 0 5108 0 1 10880
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_49
timestamp 1571791925
transform 1 0 4368 0 1 11424
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_50
timestamp 1571791925
transform 1 0 5108 0 1 13056
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_51
timestamp 1571791925
transform 1 0 4368 0 1 12512
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_52
timestamp 1571791925
transform 1 0 5108 0 1 11968
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_53
timestamp 1571791925
transform 1 0 4368 0 1 13600
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_54
timestamp 1571791925
transform 1 0 5108 0 1 15232
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_55
timestamp 1571791925
transform 1 0 4368 0 1 15776
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_56
timestamp 1571791925
transform 1 0 4368 0 1 14688
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_57
timestamp 1571791925
transform 1 0 5108 0 1 14144
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_58
timestamp 1571791925
transform 1 0 5108 0 1 16320
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_59
timestamp 1571791925
transform 1 0 4368 0 1 16864
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_60
timestamp 1571791925
transform 1 0 5108 0 1 17408
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_61
timestamp 1571791925
transform 1 0 4368 0 1 17952
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_62
timestamp 1571791925
transform 1 0 4368 0 1 19040
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_63
timestamp 1571791925
transform 1 0 5108 0 1 18496
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_64
timestamp 1571791925
transform 1 0 16368 0 1 12512
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_65
timestamp 1571791925
transform 1 0 17108 0 1 10880
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_66
timestamp 1571791925
transform 1 0 17108 0 1 11968
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_67
timestamp 1571791925
transform 1 0 16368 0 1 11424
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_68
timestamp 1571791925
transform 1 0 17108 0 1 13056
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_69
timestamp 1571791925
transform 1 0 16368 0 1 15776
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_70
timestamp 1571791925
transform 1 0 17108 0 1 14144
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_71
timestamp 1571791925
transform 1 0 16368 0 1 13600
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_72
timestamp 1571791925
transform 1 0 17108 0 1 15232
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_73
timestamp 1571791925
transform 1 0 16368 0 1 14688
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_74
timestamp 1571791925
transform 1 0 10368 0 1 12512
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_75
timestamp 1571791925
transform 1 0 11108 0 1 10880
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_76
timestamp 1571791925
transform 1 0 10368 0 1 11424
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_77
timestamp 1571791925
transform 1 0 11108 0 1 11968
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_78
timestamp 1571791925
transform 1 0 11108 0 1 13056
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_79
timestamp 1571791925
transform 1 0 11108 0 1 14144
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_80
timestamp 1571791925
transform 1 0 10368 0 1 13600
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_81
timestamp 1571791925
transform 1 0 10368 0 1 14688
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_82
timestamp 1571791925
transform 1 0 10368 0 1 15776
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_83
timestamp 1571791925
transform 1 0 11108 0 1 15232
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_84
timestamp 1571791925
transform 1 0 10368 0 1 16864
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_85
timestamp 1571791925
transform 1 0 10368 0 1 17952
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_86
timestamp 1571791925
transform 1 0 10368 0 1 19040
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_87
timestamp 1571791925
transform 1 0 11108 0 1 18496
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_88
timestamp 1571791925
transform 1 0 11108 0 1 17408
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_89
timestamp 1571791925
transform 1 0 11108 0 1 16320
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_90
timestamp 1571791925
transform 1 0 16368 0 1 16864
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_91
timestamp 1571791925
transform 1 0 16368 0 1 17952
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_92
timestamp 1571791925
transform 1 0 16368 0 1 19040
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_93
timestamp 1571791925
transform 1 0 17108 0 1 18496
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_94
timestamp 1571791925
transform 1 0 17108 0 1 16320
box -192 -48 192 48
use VIA_via2_3_2000_480_1_6_320_320  VIA_via2_3_2000_480_1_6_320_320_95
timestamp 1571791925
transform 1 0 17108 0 1 17408
box -192 -48 192 48
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_0
timestamp 1571791925
transform 1 0 16368 0 1 4896
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_1
timestamp 1571791925
transform 1 0 16368 0 1 2720
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_2
timestamp 1571791925
transform 1 0 16368 0 1 3808
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_3
timestamp 1571791925
transform 1 0 17108 0 1 3264
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_4
timestamp 1571791925
transform 1 0 17108 0 1 4352
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_5
timestamp 1571791925
transform 1 0 17108 0 1 2176
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_6
timestamp 1571791925
transform 1 0 11108 0 1 2176
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_7
timestamp 1571791925
transform 1 0 10368 0 1 2720
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_8
timestamp 1571791925
transform 1 0 10368 0 1 4896
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_9
timestamp 1571791925
transform 1 0 11108 0 1 3264
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_10
timestamp 1571791925
transform 1 0 11108 0 1 4352
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_11
timestamp 1571791925
transform 1 0 10368 0 1 3808
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_12
timestamp 1571791925
transform 1 0 11108 0 1 7616
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_13
timestamp 1571791925
transform 1 0 11108 0 1 5440
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_14
timestamp 1571791925
transform 1 0 11108 0 1 6528
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_15
timestamp 1571791925
transform 1 0 10368 0 1 5984
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_16
timestamp 1571791925
transform 1 0 10368 0 1 7072
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_17
timestamp 1571791925
transform 1 0 10368 0 1 10336
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_18
timestamp 1571791925
transform 1 0 10368 0 1 9248
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_19
timestamp 1571791925
transform 1 0 10368 0 1 8160
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_20
timestamp 1571791925
transform 1 0 11108 0 1 8704
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_21
timestamp 1571791925
transform 1 0 11108 0 1 9792
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_22
timestamp 1571791925
transform 1 0 16368 0 1 5984
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_23
timestamp 1571791925
transform 1 0 17108 0 1 7616
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_24
timestamp 1571791925
transform 1 0 16368 0 1 7072
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_25
timestamp 1571791925
transform 1 0 17108 0 1 5440
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_26
timestamp 1571791925
transform 1 0 17108 0 1 6528
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_27
timestamp 1571791925
transform 1 0 17108 0 1 8704
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_28
timestamp 1571791925
transform 1 0 17108 0 1 9792
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_29
timestamp 1571791925
transform 1 0 16368 0 1 10336
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_30
timestamp 1571791925
transform 1 0 16368 0 1 9248
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_31
timestamp 1571791925
transform 1 0 16368 0 1 8160
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_32
timestamp 1571791925
transform 1 0 5108 0 1 2176
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_33
timestamp 1571791925
transform 1 0 4368 0 1 4896
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_34
timestamp 1571791925
transform 1 0 4368 0 1 3808
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_35
timestamp 1571791925
transform 1 0 5108 0 1 4352
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_36
timestamp 1571791925
transform 1 0 4368 0 1 2720
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_37
timestamp 1571791925
transform 1 0 5108 0 1 3264
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_38
timestamp 1571791925
transform 1 0 5108 0 1 5440
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_39
timestamp 1571791925
transform 1 0 5108 0 1 6528
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_40
timestamp 1571791925
transform 1 0 5108 0 1 7616
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_41
timestamp 1571791925
transform 1 0 4368 0 1 5984
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_42
timestamp 1571791925
transform 1 0 4368 0 1 7072
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_43
timestamp 1571791925
transform 1 0 4368 0 1 9248
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_44
timestamp 1571791925
transform 1 0 4368 0 1 10336
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_45
timestamp 1571791925
transform 1 0 4368 0 1 8160
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_46
timestamp 1571791925
transform 1 0 5108 0 1 9792
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_47
timestamp 1571791925
transform 1 0 5108 0 1 8704
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_48
timestamp 1571791925
transform 1 0 4368 0 1 11424
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_49
timestamp 1571791925
transform 1 0 5108 0 1 10880
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_50
timestamp 1571791925
transform 1 0 5108 0 1 13056
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_51
timestamp 1571791925
transform 1 0 4368 0 1 12512
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_52
timestamp 1571791925
transform 1 0 5108 0 1 11968
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_53
timestamp 1571791925
transform 1 0 5108 0 1 14144
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_54
timestamp 1571791925
transform 1 0 4368 0 1 13600
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_55
timestamp 1571791925
transform 1 0 4368 0 1 15776
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_56
timestamp 1571791925
transform 1 0 4368 0 1 14688
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_57
timestamp 1571791925
transform 1 0 5108 0 1 15232
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_58
timestamp 1571791925
transform 1 0 4368 0 1 17952
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_59
timestamp 1571791925
transform 1 0 5108 0 1 18496
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_60
timestamp 1571791925
transform 1 0 4368 0 1 16864
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_61
timestamp 1571791925
transform 1 0 5108 0 1 17408
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_62
timestamp 1571791925
transform 1 0 5108 0 1 16320
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_63
timestamp 1571791925
transform 1 0 4368 0 1 19040
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_64
timestamp 1571791925
transform 1 0 17108 0 1 10880
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_65
timestamp 1571791925
transform 1 0 17108 0 1 11968
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_66
timestamp 1571791925
transform 1 0 16368 0 1 12512
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_67
timestamp 1571791925
transform 1 0 17108 0 1 13056
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_68
timestamp 1571791925
transform 1 0 16368 0 1 11424
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_69
timestamp 1571791925
transform 1 0 17108 0 1 14144
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_70
timestamp 1571791925
transform 1 0 17108 0 1 15232
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_71
timestamp 1571791925
transform 1 0 16368 0 1 14688
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_72
timestamp 1571791925
transform 1 0 16368 0 1 13600
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_73
timestamp 1571791925
transform 1 0 16368 0 1 15776
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_74
timestamp 1571791925
transform 1 0 11108 0 1 10880
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_75
timestamp 1571791925
transform 1 0 11108 0 1 11968
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_76
timestamp 1571791925
transform 1 0 11108 0 1 13056
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_77
timestamp 1571791925
transform 1 0 10368 0 1 12512
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_78
timestamp 1571791925
transform 1 0 10368 0 1 11424
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_79
timestamp 1571791925
transform 1 0 10368 0 1 14688
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_80
timestamp 1571791925
transform 1 0 11108 0 1 14144
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_81
timestamp 1571791925
transform 1 0 10368 0 1 15776
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_82
timestamp 1571791925
transform 1 0 10368 0 1 13600
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_83
timestamp 1571791925
transform 1 0 11108 0 1 15232
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_84
timestamp 1571791925
transform 1 0 11108 0 1 17408
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_85
timestamp 1571791925
transform 1 0 11108 0 1 18496
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_86
timestamp 1571791925
transform 1 0 11108 0 1 16320
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_87
timestamp 1571791925
transform 1 0 10368 0 1 17952
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_88
timestamp 1571791925
transform 1 0 10368 0 1 19040
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_89
timestamp 1571791925
transform 1 0 10368 0 1 16864
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_90
timestamp 1571791925
transform 1 0 16368 0 1 16864
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_91
timestamp 1571791925
transform 1 0 16368 0 1 19040
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_92
timestamp 1571791925
transform 1 0 16368 0 1 17952
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_93
timestamp 1571791925
transform 1 0 17108 0 1 16320
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_94
timestamp 1571791925
transform 1 0 17108 0 1 18496
box -193 -37 193 37
use VIA_via3_4_2000_480_1_5_400_400  VIA_via3_4_2000_480_1_5_400_400_95
timestamp 1571791925
transform 1 0 17108 0 1 17408
box -193 -37 193 37
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_0
timestamp 1571791925
transform 1 0 17108 0 1 3264
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_1
timestamp 1571791925
transform 1 0 17108 0 1 2176
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_2
timestamp 1571791925
transform 1 0 16368 0 1 2720
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_3
timestamp 1571791925
transform 1 0 16368 0 1 3808
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_4
timestamp 1571791925
transform 1 0 17108 0 1 4352
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_5
timestamp 1571791925
transform 1 0 16368 0 1 4896
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_6
timestamp 1571791925
transform 1 0 11108 0 1 2176
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_7
timestamp 1571791925
transform 1 0 11108 0 1 4352
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_8
timestamp 1571791925
transform 1 0 11108 0 1 3264
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_9
timestamp 1571791925
transform 1 0 10368 0 1 3808
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_10
timestamp 1571791925
transform 1 0 10368 0 1 2720
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_11
timestamp 1571791925
transform 1 0 10368 0 1 4896
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_12
timestamp 1571791925
transform 1 0 11108 0 1 7616
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_13
timestamp 1571791925
transform 1 0 11108 0 1 5440
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_14
timestamp 1571791925
transform 1 0 10368 0 1 7072
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_15
timestamp 1571791925
transform 1 0 11108 0 1 6528
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_16
timestamp 1571791925
transform 1 0 10368 0 1 5984
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_17
timestamp 1571791925
transform 1 0 10368 0 1 9248
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_18
timestamp 1571791925
transform 1 0 10368 0 1 8160
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_19
timestamp 1571791925
transform 1 0 10368 0 1 10336
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_20
timestamp 1571791925
transform 1 0 11108 0 1 8704
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_21
timestamp 1571791925
transform 1 0 11108 0 1 9792
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_22
timestamp 1571791925
transform 1 0 17108 0 1 6528
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_23
timestamp 1571791925
transform 1 0 16368 0 1 5984
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_24
timestamp 1571791925
transform 1 0 17108 0 1 7616
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_25
timestamp 1571791925
transform 1 0 17108 0 1 5440
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_26
timestamp 1571791925
transform 1 0 16368 0 1 7072
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_27
timestamp 1571791925
transform 1 0 16368 0 1 10336
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_28
timestamp 1571791925
transform 1 0 16368 0 1 8160
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_29
timestamp 1571791925
transform 1 0 16368 0 1 9248
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_30
timestamp 1571791925
transform 1 0 17108 0 1 8704
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_31
timestamp 1571791925
transform 1 0 17108 0 1 9792
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_32
timestamp 1571791925
transform 1 0 5108 0 1 2176
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_33
timestamp 1571791925
transform 1 0 4368 0 1 4896
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_34
timestamp 1571791925
transform 1 0 5108 0 1 3264
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_35
timestamp 1571791925
transform 1 0 5108 0 1 4352
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_36
timestamp 1571791925
transform 1 0 4368 0 1 2720
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_37
timestamp 1571791925
transform 1 0 4368 0 1 3808
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_38
timestamp 1571791925
transform 1 0 4368 0 1 7072
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_39
timestamp 1571791925
transform 1 0 5108 0 1 7616
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_40
timestamp 1571791925
transform 1 0 5108 0 1 5440
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_41
timestamp 1571791925
transform 1 0 5108 0 1 6528
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_42
timestamp 1571791925
transform 1 0 4368 0 1 5984
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_43
timestamp 1571791925
transform 1 0 4368 0 1 9248
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_44
timestamp 1571791925
transform 1 0 4368 0 1 10336
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_45
timestamp 1571791925
transform 1 0 5108 0 1 8704
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_46
timestamp 1571791925
transform 1 0 5108 0 1 9792
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_47
timestamp 1571791925
transform 1 0 4368 0 1 8160
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_48
timestamp 1571791925
transform 1 0 5108 0 1 11968
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_49
timestamp 1571791925
transform 1 0 4368 0 1 12512
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_50
timestamp 1571791925
transform 1 0 5108 0 1 13056
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_51
timestamp 1571791925
transform 1 0 5108 0 1 10880
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_52
timestamp 1571791925
transform 1 0 4368 0 1 11424
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_53
timestamp 1571791925
transform 1 0 4368 0 1 13600
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_54
timestamp 1571791925
transform 1 0 4368 0 1 14688
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_55
timestamp 1571791925
transform 1 0 4368 0 1 15776
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_56
timestamp 1571791925
transform 1 0 5108 0 1 15232
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_57
timestamp 1571791925
transform 1 0 5108 0 1 14144
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_58
timestamp 1571791925
transform 1 0 5108 0 1 16320
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_59
timestamp 1571791925
transform 1 0 5108 0 1 17408
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_60
timestamp 1571791925
transform 1 0 4368 0 1 17952
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_61
timestamp 1571791925
transform 1 0 4368 0 1 16864
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_62
timestamp 1571791925
transform 1 0 5108 0 1 18496
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_63
timestamp 1571791925
transform 1 0 4368 0 1 19040
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_64
timestamp 1571791925
transform 1 0 17108 0 1 10880
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_65
timestamp 1571791925
transform 1 0 17108 0 1 13056
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_66
timestamp 1571791925
transform 1 0 17108 0 1 11968
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_67
timestamp 1571791925
transform 1 0 16368 0 1 11424
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_68
timestamp 1571791925
transform 1 0 16368 0 1 12512
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_69
timestamp 1571791925
transform 1 0 16368 0 1 14688
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_70
timestamp 1571791925
transform 1 0 17108 0 1 14144
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_71
timestamp 1571791925
transform 1 0 16368 0 1 15776
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_72
timestamp 1571791925
transform 1 0 16368 0 1 13600
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_73
timestamp 1571791925
transform 1 0 17108 0 1 15232
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_74
timestamp 1571791925
transform 1 0 11108 0 1 13056
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_75
timestamp 1571791925
transform 1 0 11108 0 1 11968
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_76
timestamp 1571791925
transform 1 0 11108 0 1 10880
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_77
timestamp 1571791925
transform 1 0 10368 0 1 11424
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_78
timestamp 1571791925
transform 1 0 10368 0 1 12512
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_79
timestamp 1571791925
transform 1 0 10368 0 1 14688
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_80
timestamp 1571791925
transform 1 0 11108 0 1 14144
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_81
timestamp 1571791925
transform 1 0 11108 0 1 15232
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_82
timestamp 1571791925
transform 1 0 10368 0 1 15776
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_83
timestamp 1571791925
transform 1 0 10368 0 1 13600
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_84
timestamp 1571791925
transform 1 0 10368 0 1 17952
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_85
timestamp 1571791925
transform 1 0 10368 0 1 19040
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_86
timestamp 1571791925
transform 1 0 10368 0 1 16864
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_87
timestamp 1571791925
transform 1 0 11108 0 1 18496
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_88
timestamp 1571791925
transform 1 0 11108 0 1 17408
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_89
timestamp 1571791925
transform 1 0 11108 0 1 16320
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_90
timestamp 1571791925
transform 1 0 16368 0 1 19040
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_91
timestamp 1571791925
transform 1 0 16368 0 1 16864
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_92
timestamp 1571791925
transform 1 0 16368 0 1 17952
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_93
timestamp 1571791925
transform 1 0 17108 0 1 16320
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_94
timestamp 1571791925
transform 1 0 17108 0 1 18496
box -200 -33 200 33
use VIA_via4_5_2000_480_1_5_400_400  VIA_via4_5_2000_480_1_5_400_400_95
timestamp 1571791925
transform 1 0 17108 0 1 17408
box -200 -33 200 33
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_0
timestamp 1571791925
transform 1 0 11108 0 1 6246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_1
timestamp 1571791925
transform 1 0 17108 0 1 6246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_2
timestamp 1571791925
transform 1 0 10368 0 1 5506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_3
timestamp 1571791925
transform 1 0 16368 0 1 5506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_4
timestamp 1571791925
transform 1 0 5108 0 1 6246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_5
timestamp 1571791925
transform 1 0 4368 0 1 5506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_6
timestamp 1571791925
transform 1 0 4368 0 1 11506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_7
timestamp 1571791925
transform 1 0 5108 0 1 12246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_8
timestamp 1571791925
transform 1 0 5108 0 1 18246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_9
timestamp 1571791925
transform 1 0 4368 0 1 17506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_10
timestamp 1571791925
transform 1 0 17108 0 1 12246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_11
timestamp 1571791925
transform 1 0 16368 0 1 11506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_12
timestamp 1571791925
transform 1 0 10368 0 1 11506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_13
timestamp 1571791925
transform 1 0 11108 0 1 12246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_14
timestamp 1571791925
transform 1 0 11108 0 1 18246
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_15
timestamp 1571791925
transform 1 0 10368 0 1 17506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_16
timestamp 1571791925
transform 1 0 16368 0 1 17506
box -200 -200 200 200
use VIA_via5_6_2000_2000_1_1_1600_1600  VIA_via5_6_2000_2000_1_1_1600_1600_17
timestamp 1571791925
transform 1 0 17108 0 1 18246
box -200 -200 200 200
<< labels >>
rlabel metal3 s 0 21088 800 21208 4 clk
port 2 nsew
rlabel metal3 s 0 20408 800 20528 4 p
port 3 nsew
rlabel metal3 s 0 19728 800 19848 4 rst
port 4 nsew
rlabel metal3 s 0 19048 800 19168 4 x[0]
port 5 nsew
rlabel metal3 s 0 18368 800 18488 4 x[10]
port 6 nsew
rlabel metal3 s 0 17688 800 17808 4 x[11]
port 7 nsew
rlabel metal3 s 0 17008 800 17128 4 x[12]
port 8 nsew
rlabel metal3 s 0 16328 800 16448 4 x[13]
port 9 nsew
rlabel metal3 s 0 15648 800 15768 4 x[14]
port 10 nsew
rlabel metal3 s 0 14968 800 15088 4 x[15]
port 11 nsew
rlabel metal3 s 0 14288 800 14408 4 x[16]
port 12 nsew
rlabel metal3 s 0 13608 800 13728 4 x[17]
port 13 nsew
rlabel metal3 s 0 12928 800 13048 4 x[18]
port 14 nsew
rlabel metal3 s 0 12248 800 12368 4 x[19]
port 15 nsew
rlabel metal3 s 0 11568 800 11688 4 x[1]
port 16 nsew
rlabel metal3 s 0 10888 800 11008 4 x[20]
port 17 nsew
rlabel metal3 s 0 10208 800 10328 4 x[21]
port 18 nsew
rlabel metal3 s 0 9528 800 9648 4 x[22]
port 19 nsew
rlabel metal3 s 0 8848 800 8968 4 x[23]
port 20 nsew
rlabel metal3 s 0 8168 800 8288 4 x[24]
port 21 nsew
rlabel metal3 s 0 7488 800 7608 4 x[25]
port 22 nsew
rlabel metal3 s 0 6808 800 6928 4 x[26]
port 23 nsew
rlabel metal3 s 0 6128 800 6248 4 x[27]
port 24 nsew
rlabel metal3 s 0 5448 800 5568 4 x[28]
port 25 nsew
rlabel metal3 s 0 4768 800 4888 4 x[29]
port 26 nsew
rlabel metal3 s 0 4088 800 4208 4 x[2]
port 27 nsew
rlabel metal3 s 0 3408 800 3528 4 x[30]
port 28 nsew
rlabel metal3 s 0 2728 800 2848 4 x[31]
port 29 nsew
rlabel metal3 s 0 2048 800 2168 4 x[3]
port 30 nsew
rlabel metal3 s 0 1368 800 1488 4 x[4]
port 31 nsew
rlabel metal3 s 0 688 800 808 4 x[5]
port 32 nsew
rlabel metal3 s 0 8 800 128 4 x[6]
port 33 nsew
rlabel metal3 s 18507 9528 19307 9648 4 x[7]
port 34 nsew
rlabel metal3 s 18507 10888 19307 11008 4 x[8]
port 35 nsew
rlabel metal3 s 18507 10208 19307 10328 4 x[9]
port 36 nsew
rlabel metal3 s 18507 11568 19307 11688 4 y
port 37 nsew
rlabel metal4 s 4908 2128 5308 19088 4 VGND
port 39 nsew
rlabel metal4 s 4168 2128 4568 19088 4 VPWR
port 40 nsew
rlabel metal5 s 1056 6046 18172 6446 4 VGND
port 39 nsew
rlabel metal5 s 1056 5306 18172 5706 4 VPWR
port 40 nsew
<< properties >>
string FIXED_BBOX 0 0 19307 21451
string path 5.280 27.530 90.860 27.530 
<< end >>
